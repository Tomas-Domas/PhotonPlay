module rom_dev #(
    parameter LUT_SIZE = 4096
)
(
    input clk,
    input we,
    input [$clog2(LUT_SIZE)-1:0] addr,
    input [11:0] di,
    output [11:0] dout
);

    reg [11:0] rom [LUT_SIZE-1:0];
    reg [11:0] dout;

    initial begin
        rom[0] = 12'd4095;
        rom[1] = 12'd4093;
        rom[2] = 12'd4085;
        rom[3] = 12'd4073;
        rom[4] = 12'd4056;
        rom[5] = 12'd4034;
        rom[6] = 12'd4007;
        rom[7] = 12'd3975;
        rom[8] = 12'd3939;
        rom[9] = 12'd3898;
        rom[10] = 12'd3853;
        rom[11] = 12'd3804;
        rom[12] = 12'd3750;
        rom[13] = 12'd3692;
        rom[14] = 12'd3630;
        rom[15] = 12'd3565;
        rom[16] = 12'd3495;
        rom[17] = 12'd3423;
        rom[18] = 12'd3346;
        rom[19] = 12'd3267;
        rom[20] = 12'd3185;
        rom[21] = 12'd3100;
        rom[22] = 12'd3013;
        rom[23] = 12'd2923;
        rom[24] = 12'd2831;
        rom[25] = 12'd2737;
        rom[26] = 12'd2642;
        rom[27] = 12'd2545;
        rom[28] = 12'd2447;
        rom[29] = 12'd2348;
        rom[30] = 12'd2248;
        rom[31] = 12'd2148;
        rom[32] = 12'd2048;
        rom[33] = 12'd1947;
        rom[34] = 12'd1847;
        rom[35] = 12'd1747;
        rom[36] = 12'd1648;
        rom[37] = 12'd1550;
        rom[38] = 12'd1453;
        rom[39] = 12'd1358;
        rom[40] = 12'd1264;
        rom[41] = 12'd1172;
        rom[42] = 12'd1082;
        rom[43] = 12'd995;
        rom[44] = 12'd910;
        rom[45] = 12'd828;
        rom[46] = 12'd749;
        rom[47] = 12'd672;
        rom[48] = 12'd600;
        rom[49] = 12'd530;
        rom[50] = 12'd465;
        rom[51] = 12'd403;
        rom[52] = 12'd345;
        rom[53] = 12'd291;
        rom[54] = 12'd242;
        rom[55] = 12'd197;
        rom[56] = 12'd156;
        rom[57] = 12'd120;
        rom[58] = 12'd88;
        rom[59] = 12'd61;
        rom[60] = 12'd39;
        rom[61] = 12'd22;
        rom[62] = 12'd10;
        rom[63] = 12'd2;
        rom[64] = 12'd0;
        rom[65] = 12'd2;
        rom[66] = 12'd10;
        rom[67] = 12'd22;
        rom[68] = 12'd39;
        rom[69] = 12'd61;
        rom[70] = 12'd88;
        rom[71] = 12'd120;
        rom[72] = 12'd156;
        rom[73] = 12'd197;
        rom[74] = 12'd242;
        rom[75] = 12'd291;
        rom[76] = 12'd345;
        rom[77] = 12'd403;
        rom[78] = 12'd465;
        rom[79] = 12'd530;
        rom[80] = 12'd600;
        rom[81] = 12'd672;
        rom[82] = 12'd749;
        rom[83] = 12'd828;
        rom[84] = 12'd910;
        rom[85] = 12'd995;
        rom[86] = 12'd1082;
        rom[87] = 12'd1172;
        rom[88] = 12'd1264;
        rom[89] = 12'd1358;
        rom[90] = 12'd1453;
        rom[91] = 12'd1550;
        rom[92] = 12'd1648;
        rom[93] = 12'd1747;
        rom[94] = 12'd1847;
        rom[95] = 12'd1947;
        rom[96] = 12'd2047;
        rom[97] = 12'd2148;
        rom[98] = 12'd2248;
        rom[99] = 12'd2348;
        rom[100] = 12'd2447;
        rom[101] = 12'd2545;
        rom[102] = 12'd2642;
        rom[103] = 12'd2737;
        rom[104] = 12'd2831;
        rom[105] = 12'd2923;
        rom[106] = 12'd3013;
        rom[107] = 12'd3100;
        rom[108] = 12'd3185;
        rom[109] = 12'd3267;
        rom[110] = 12'd3346;
        rom[111] = 12'd3423;
        rom[112] = 12'd3495;
        rom[113] = 12'd3565;
        rom[114] = 12'd3630;
        rom[115] = 12'd3692;
        rom[116] = 12'd3750;
        rom[117] = 12'd3804;
        rom[118] = 12'd3853;
        rom[119] = 12'd3898;
        rom[120] = 12'd3939;
        rom[121] = 12'd3975;
        rom[122] = 12'd4007;
        rom[123] = 12'd4034;
        rom[124] = 12'd4056;
        rom[125] = 12'd4073;
        rom[126] = 12'd4085;
        rom[127] = 12'd4093;
    end

    always @(posedge clk) begin
        if (we) rom[addr] <= di;
        dout <= rom[addr];
    end

endmodule