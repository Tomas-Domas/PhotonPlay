module rom_dev #(
    localparam LUT_SIZE = 4096
)
(
    input clk,
    input we,
    input [$clog2(LUT_SIZE)-1:0] addr,
    input [11:0] di,
    output [11:0] dout
);

    reg [11:0] rom [LUT_SIZE-1:0];
    reg [11:0] dout;

    initial begin
        rom[0] = 12'd0;
        rom[1] = 12'd1;
        rom[2] = 12'd2;
        rom[3] = 12'd3;
        rom[4] = 12'd4;
        rom[5] = 12'd5;
        rom[6] = 12'd6;
        rom[7] = 12'd7;
        rom[8] = 12'd8;
        rom[9] = 12'd9;
        rom[10] = 12'd10;
        rom[11] = 12'd11;
        rom[12] = 12'd12;
        rom[13] = 12'd13;
        rom[14] = 12'd14;
        rom[15] = 12'd15;
        rom[16] = 12'd16;
        rom[17] = 12'd17;
        rom[18] = 12'd18;
        rom[19] = 12'd19;
        rom[20] = 12'd20;
        rom[21] = 12'd21;
        rom[22] = 12'd22;
        rom[23] = 12'd23;
        rom[24] = 12'd24;
        rom[25] = 12'd25;
        rom[26] = 12'd26;
        rom[27] = 12'd27;
        rom[28] = 12'd28;
        rom[29] = 12'd29;
        rom[30] = 12'd30;
        rom[31] = 12'd31;
        rom[32] = 12'd32;
        rom[33] = 12'd33;
        rom[34] = 12'd34;
        rom[35] = 12'd35;
        rom[36] = 12'd36;
        rom[37] = 12'd37;
        rom[38] = 12'd38;
        rom[39] = 12'd39;
        rom[40] = 12'd40;
        rom[41] = 12'd41;
        rom[42] = 12'd42;
        rom[43] = 12'd43;
        rom[44] = 12'd44;
        rom[45] = 12'd45;
        rom[46] = 12'd46;
        rom[47] = 12'd47;
        rom[48] = 12'd48;
        rom[49] = 12'd49;
        rom[50] = 12'd50;
        rom[51] = 12'd51;
        rom[52] = 12'd52;
        rom[53] = 12'd53;
        rom[54] = 12'd54;
        rom[55] = 12'd55;
        rom[56] = 12'd56;
        rom[57] = 12'd57;
        rom[58] = 12'd58;
        rom[59] = 12'd59;
        rom[60] = 12'd60;
        rom[61] = 12'd61;
        rom[62] = 12'd62;
        rom[63] = 12'd63;
        rom[64] = 12'd64;
        rom[65] = 12'd65;
        rom[66] = 12'd66;
        rom[67] = 12'd67;
        rom[68] = 12'd68;
        rom[69] = 12'd69;
        rom[70] = 12'd70;
        rom[71] = 12'd71;
        rom[72] = 12'd72;
        rom[73] = 12'd73;
        rom[74] = 12'd74;
        rom[75] = 12'd75;
        rom[76] = 12'd76;
        rom[77] = 12'd77;
        rom[78] = 12'd78;
        rom[79] = 12'd79;
        rom[80] = 12'd80;
        rom[81] = 12'd81;
        rom[82] = 12'd82;
        rom[83] = 12'd83;
        rom[84] = 12'd84;
        rom[85] = 12'd85;
        rom[86] = 12'd86;
        rom[87] = 12'd87;
        rom[88] = 12'd88;
        rom[89] = 12'd89;
        rom[90] = 12'd90;
        rom[91] = 12'd91;
        rom[92] = 12'd92;
        rom[93] = 12'd93;
        rom[94] = 12'd94;
        rom[95] = 12'd95;
        rom[96] = 12'd96;
        rom[97] = 12'd97;
        rom[98] = 12'd98;
        rom[99] = 12'd99;
        rom[100] = 12'd100;
        rom[101] = 12'd101;
        rom[102] = 12'd102;
        rom[103] = 12'd103;
        rom[104] = 12'd104;
        rom[105] = 12'd105;
        rom[106] = 12'd106;
        rom[107] = 12'd107;
        rom[108] = 12'd108;
        rom[109] = 12'd109;
        rom[110] = 12'd110;
        rom[111] = 12'd111;
        rom[112] = 12'd112;
        rom[113] = 12'd113;
        rom[114] = 12'd114;
        rom[115] = 12'd115;
        rom[116] = 12'd116;
        rom[117] = 12'd117;
        rom[118] = 12'd118;
        rom[119] = 12'd119;
        rom[120] = 12'd120;
        rom[121] = 12'd121;
        rom[122] = 12'd122;
        rom[123] = 12'd123;
        rom[124] = 12'd124;
        rom[125] = 12'd125;
        rom[126] = 12'd126;
        rom[127] = 12'd127;
        rom[128] = 12'd128;
        rom[129] = 12'd129;
        rom[130] = 12'd130;
        rom[131] = 12'd131;
        rom[132] = 12'd132;
        rom[133] = 12'd133;
        rom[134] = 12'd134;
        rom[135] = 12'd135;
        rom[136] = 12'd136;
        rom[137] = 12'd137;
        rom[138] = 12'd138;
        rom[139] = 12'd139;
        rom[140] = 12'd140;
        rom[141] = 12'd141;
        rom[142] = 12'd142;
        rom[143] = 12'd143;
        rom[144] = 12'd144;
        rom[145] = 12'd145;
        rom[146] = 12'd146;
        rom[147] = 12'd147;
        rom[148] = 12'd148;
        rom[149] = 12'd149;
        rom[150] = 12'd150;
        rom[151] = 12'd151;
        rom[152] = 12'd152;
        rom[153] = 12'd153;
        rom[154] = 12'd154;
        rom[155] = 12'd155;
        rom[156] = 12'd156;
        rom[157] = 12'd157;
        rom[158] = 12'd158;
        rom[159] = 12'd159;
        rom[160] = 12'd160;
        rom[161] = 12'd161;
        rom[162] = 12'd162;
        rom[163] = 12'd163;
        rom[164] = 12'd164;
        rom[165] = 12'd165;
        rom[166] = 12'd166;
        rom[167] = 12'd167;
        rom[168] = 12'd168;
        rom[169] = 12'd169;
        rom[170] = 12'd170;
        rom[171] = 12'd171;
        rom[172] = 12'd172;
        rom[173] = 12'd173;
        rom[174] = 12'd174;
        rom[175] = 12'd175;
        rom[176] = 12'd176;
        rom[177] = 12'd177;
        rom[178] = 12'd178;
        rom[179] = 12'd179;
        rom[180] = 12'd180;
        rom[181] = 12'd181;
        rom[182] = 12'd182;
        rom[183] = 12'd183;
        rom[184] = 12'd184;
        rom[185] = 12'd185;
        rom[186] = 12'd186;
        rom[187] = 12'd187;
        rom[188] = 12'd188;
        rom[189] = 12'd189;
        rom[190] = 12'd190;
        rom[191] = 12'd191;
        rom[192] = 12'd192;
        rom[193] = 12'd193;
        rom[194] = 12'd194;
        rom[195] = 12'd195;
        rom[196] = 12'd196;
        rom[197] = 12'd197;
        rom[198] = 12'd198;
        rom[199] = 12'd199;
        rom[200] = 12'd200;
        rom[201] = 12'd201;
        rom[202] = 12'd202;
        rom[203] = 12'd203;
        rom[204] = 12'd204;
        rom[205] = 12'd205;
        rom[206] = 12'd206;
        rom[207] = 12'd207;
        rom[208] = 12'd208;
        rom[209] = 12'd209;
        rom[210] = 12'd210;
        rom[211] = 12'd211;
        rom[212] = 12'd212;
        rom[213] = 12'd213;
        rom[214] = 12'd214;
        rom[215] = 12'd215;
        rom[216] = 12'd216;
        rom[217] = 12'd217;
        rom[218] = 12'd218;
        rom[219] = 12'd219;
        rom[220] = 12'd220;
        rom[221] = 12'd221;
        rom[222] = 12'd222;
        rom[223] = 12'd223;
        rom[224] = 12'd224;
        rom[225] = 12'd225;
        rom[226] = 12'd226;
        rom[227] = 12'd227;
        rom[228] = 12'd228;
        rom[229] = 12'd229;
        rom[230] = 12'd230;
        rom[231] = 12'd231;
        rom[232] = 12'd232;
        rom[233] = 12'd233;
        rom[234] = 12'd234;
        rom[235] = 12'd235;
        rom[236] = 12'd236;
        rom[237] = 12'd237;
        rom[238] = 12'd238;
        rom[239] = 12'd239;
        rom[240] = 12'd240;
        rom[241] = 12'd241;
        rom[242] = 12'd242;
        rom[243] = 12'd243;
        rom[244] = 12'd244;
        rom[245] = 12'd245;
        rom[246] = 12'd246;
        rom[247] = 12'd247;
        rom[248] = 12'd248;
        rom[249] = 12'd249;
        rom[250] = 12'd250;
        rom[251] = 12'd251;
        rom[252] = 12'd252;
        rom[253] = 12'd253;
        rom[254] = 12'd254;
        rom[255] = 12'd255;
        rom[256] = 12'd256;
        rom[257] = 12'd257;
        rom[258] = 12'd258;
        rom[259] = 12'd259;
        rom[260] = 12'd260;
        rom[261] = 12'd261;
        rom[262] = 12'd262;
        rom[263] = 12'd263;
        rom[264] = 12'd264;
        rom[265] = 12'd265;
        rom[266] = 12'd266;
        rom[267] = 12'd267;
        rom[268] = 12'd268;
        rom[269] = 12'd269;
        rom[270] = 12'd270;
        rom[271] = 12'd271;
        rom[272] = 12'd272;
        rom[273] = 12'd273;
        rom[274] = 12'd274;
        rom[275] = 12'd275;
        rom[276] = 12'd276;
        rom[277] = 12'd277;
        rom[278] = 12'd278;
        rom[279] = 12'd279;
        rom[280] = 12'd280;
        rom[281] = 12'd281;
        rom[282] = 12'd282;
        rom[283] = 12'd283;
        rom[284] = 12'd284;
        rom[285] = 12'd285;
        rom[286] = 12'd286;
        rom[287] = 12'd287;
        rom[288] = 12'd288;
        rom[289] = 12'd289;
        rom[290] = 12'd290;
        rom[291] = 12'd291;
        rom[292] = 12'd292;
        rom[293] = 12'd293;
        rom[294] = 12'd294;
        rom[295] = 12'd295;
        rom[296] = 12'd296;
        rom[297] = 12'd297;
        rom[298] = 12'd298;
        rom[299] = 12'd299;
        rom[300] = 12'd300;
        rom[301] = 12'd301;
        rom[302] = 12'd302;
        rom[303] = 12'd303;
        rom[304] = 12'd304;
        rom[305] = 12'd305;
        rom[306] = 12'd306;
        rom[307] = 12'd307;
        rom[308] = 12'd308;
        rom[309] = 12'd309;
        rom[310] = 12'd310;
        rom[311] = 12'd311;
        rom[312] = 12'd312;
        rom[313] = 12'd313;
        rom[314] = 12'd314;
        rom[315] = 12'd315;
        rom[316] = 12'd316;
        rom[317] = 12'd317;
        rom[318] = 12'd318;
        rom[319] = 12'd319;
        rom[320] = 12'd320;
        rom[321] = 12'd321;
        rom[322] = 12'd322;
        rom[323] = 12'd323;
        rom[324] = 12'd324;
        rom[325] = 12'd325;
        rom[326] = 12'd326;
        rom[327] = 12'd327;
        rom[328] = 12'd328;
        rom[329] = 12'd329;
        rom[330] = 12'd330;
        rom[331] = 12'd331;
        rom[332] = 12'd332;
        rom[333] = 12'd333;
        rom[334] = 12'd334;
        rom[335] = 12'd335;
        rom[336] = 12'd336;
        rom[337] = 12'd337;
        rom[338] = 12'd338;
        rom[339] = 12'd339;
        rom[340] = 12'd340;
        rom[341] = 12'd341;
        rom[342] = 12'd342;
        rom[343] = 12'd343;
        rom[344] = 12'd344;
        rom[345] = 12'd345;
        rom[346] = 12'd346;
        rom[347] = 12'd347;
        rom[348] = 12'd348;
        rom[349] = 12'd349;
        rom[350] = 12'd350;
        rom[351] = 12'd351;
        rom[352] = 12'd352;
        rom[353] = 12'd353;
        rom[354] = 12'd354;
        rom[355] = 12'd355;
        rom[356] = 12'd356;
        rom[357] = 12'd357;
        rom[358] = 12'd358;
        rom[359] = 12'd359;
        rom[360] = 12'd360;
        rom[361] = 12'd361;
        rom[362] = 12'd362;
        rom[363] = 12'd363;
        rom[364] = 12'd364;
        rom[365] = 12'd365;
        rom[366] = 12'd366;
        rom[367] = 12'd367;
        rom[368] = 12'd368;
        rom[369] = 12'd369;
        rom[370] = 12'd370;
        rom[371] = 12'd371;
        rom[372] = 12'd372;
        rom[373] = 12'd373;
        rom[374] = 12'd374;
        rom[375] = 12'd375;
        rom[376] = 12'd376;
        rom[377] = 12'd377;
        rom[378] = 12'd378;
        rom[379] = 12'd379;
        rom[380] = 12'd380;
        rom[381] = 12'd381;
        rom[382] = 12'd382;
        rom[383] = 12'd383;
        rom[384] = 12'd384;
        rom[385] = 12'd385;
        rom[386] = 12'd386;
        rom[387] = 12'd387;
        rom[388] = 12'd388;
        rom[389] = 12'd389;
        rom[390] = 12'd390;
        rom[391] = 12'd391;
        rom[392] = 12'd392;
        rom[393] = 12'd393;
        rom[394] = 12'd394;
        rom[395] = 12'd395;
        rom[396] = 12'd396;
        rom[397] = 12'd397;
        rom[398] = 12'd398;
        rom[399] = 12'd399;
        rom[400] = 12'd400;
        rom[401] = 12'd401;
        rom[402] = 12'd402;
        rom[403] = 12'd403;
        rom[404] = 12'd404;
        rom[405] = 12'd405;
        rom[406] = 12'd406;
        rom[407] = 12'd407;
        rom[408] = 12'd408;
        rom[409] = 12'd409;
        rom[410] = 12'd410;
        rom[411] = 12'd411;
        rom[412] = 12'd412;
        rom[413] = 12'd413;
        rom[414] = 12'd414;
        rom[415] = 12'd415;
        rom[416] = 12'd416;
        rom[417] = 12'd417;
        rom[418] = 12'd418;
        rom[419] = 12'd419;
        rom[420] = 12'd420;
        rom[421] = 12'd421;
        rom[422] = 12'd422;
        rom[423] = 12'd423;
        rom[424] = 12'd424;
        rom[425] = 12'd425;
        rom[426] = 12'd426;
        rom[427] = 12'd427;
        rom[428] = 12'd428;
        rom[429] = 12'd429;
        rom[430] = 12'd430;
        rom[431] = 12'd431;
        rom[432] = 12'd432;
        rom[433] = 12'd433;
        rom[434] = 12'd434;
        rom[435] = 12'd435;
        rom[436] = 12'd436;
        rom[437] = 12'd437;
        rom[438] = 12'd438;
        rom[439] = 12'd439;
        rom[440] = 12'd440;
        rom[441] = 12'd441;
        rom[442] = 12'd442;
        rom[443] = 12'd443;
        rom[444] = 12'd444;
        rom[445] = 12'd445;
        rom[446] = 12'd446;
        rom[447] = 12'd447;
        rom[448] = 12'd448;
        rom[449] = 12'd449;
        rom[450] = 12'd450;
        rom[451] = 12'd451;
        rom[452] = 12'd452;
        rom[453] = 12'd453;
        rom[454] = 12'd454;
        rom[455] = 12'd455;
        rom[456] = 12'd456;
        rom[457] = 12'd457;
        rom[458] = 12'd458;
        rom[459] = 12'd459;
        rom[460] = 12'd460;
        rom[461] = 12'd461;
        rom[462] = 12'd462;
        rom[463] = 12'd463;
        rom[464] = 12'd464;
        rom[465] = 12'd465;
        rom[466] = 12'd466;
        rom[467] = 12'd467;
        rom[468] = 12'd468;
        rom[469] = 12'd469;
        rom[470] = 12'd470;
        rom[471] = 12'd471;
        rom[472] = 12'd472;
        rom[473] = 12'd473;
        rom[474] = 12'd474;
        rom[475] = 12'd475;
        rom[476] = 12'd476;
        rom[477] = 12'd477;
        rom[478] = 12'd478;
        rom[479] = 12'd479;
        rom[480] = 12'd480;
        rom[481] = 12'd481;
        rom[482] = 12'd482;
        rom[483] = 12'd483;
        rom[484] = 12'd484;
        rom[485] = 12'd485;
        rom[486] = 12'd486;
        rom[487] = 12'd487;
        rom[488] = 12'd488;
        rom[489] = 12'd489;
        rom[490] = 12'd490;
        rom[491] = 12'd491;
        rom[492] = 12'd492;
        rom[493] = 12'd493;
        rom[494] = 12'd494;
        rom[495] = 12'd495;
        rom[496] = 12'd496;
        rom[497] = 12'd497;
        rom[498] = 12'd498;
        rom[499] = 12'd499;
        rom[500] = 12'd500;
        rom[501] = 12'd501;
        rom[502] = 12'd502;
        rom[503] = 12'd503;
        rom[504] = 12'd504;
        rom[505] = 12'd505;
        rom[506] = 12'd506;
        rom[507] = 12'd507;
        rom[508] = 12'd508;
        rom[509] = 12'd509;
        rom[510] = 12'd510;
        rom[511] = 12'd511;
        rom[512] = 12'd512;
        rom[513] = 12'd513;
        rom[514] = 12'd514;
        rom[515] = 12'd515;
        rom[516] = 12'd516;
        rom[517] = 12'd517;
        rom[518] = 12'd518;
        rom[519] = 12'd519;
        rom[520] = 12'd520;
        rom[521] = 12'd521;
        rom[522] = 12'd522;
        rom[523] = 12'd523;
        rom[524] = 12'd524;
        rom[525] = 12'd525;
        rom[526] = 12'd526;
        rom[527] = 12'd527;
        rom[528] = 12'd528;
        rom[529] = 12'd529;
        rom[530] = 12'd530;
        rom[531] = 12'd531;
        rom[532] = 12'd532;
        rom[533] = 12'd533;
        rom[534] = 12'd534;
        rom[535] = 12'd535;
        rom[536] = 12'd536;
        rom[537] = 12'd537;
        rom[538] = 12'd538;
        rom[539] = 12'd539;
        rom[540] = 12'd540;
        rom[541] = 12'd541;
        rom[542] = 12'd542;
        rom[543] = 12'd543;
        rom[544] = 12'd544;
        rom[545] = 12'd545;
        rom[546] = 12'd546;
        rom[547] = 12'd547;
        rom[548] = 12'd548;
        rom[549] = 12'd549;
        rom[550] = 12'd550;
        rom[551] = 12'd551;
        rom[552] = 12'd552;
        rom[553] = 12'd553;
        rom[554] = 12'd554;
        rom[555] = 12'd555;
        rom[556] = 12'd556;
        rom[557] = 12'd557;
        rom[558] = 12'd558;
        rom[559] = 12'd559;
        rom[560] = 12'd560;
        rom[561] = 12'd561;
        rom[562] = 12'd562;
        rom[563] = 12'd563;
        rom[564] = 12'd564;
        rom[565] = 12'd565;
        rom[566] = 12'd566;
        rom[567] = 12'd567;
        rom[568] = 12'd568;
        rom[569] = 12'd569;
        rom[570] = 12'd570;
        rom[571] = 12'd571;
        rom[572] = 12'd572;
        rom[573] = 12'd573;
        rom[574] = 12'd574;
        rom[575] = 12'd575;
        rom[576] = 12'd576;
        rom[577] = 12'd577;
        rom[578] = 12'd578;
        rom[579] = 12'd579;
        rom[580] = 12'd580;
        rom[581] = 12'd581;
        rom[582] = 12'd582;
        rom[583] = 12'd583;
        rom[584] = 12'd584;
        rom[585] = 12'd585;
        rom[586] = 12'd586;
        rom[587] = 12'd587;
        rom[588] = 12'd588;
        rom[589] = 12'd589;
        rom[590] = 12'd590;
        rom[591] = 12'd591;
        rom[592] = 12'd592;
        rom[593] = 12'd593;
        rom[594] = 12'd594;
        rom[595] = 12'd595;
        rom[596] = 12'd596;
        rom[597] = 12'd597;
        rom[598] = 12'd598;
        rom[599] = 12'd599;
        rom[600] = 12'd600;
        rom[601] = 12'd601;
        rom[602] = 12'd602;
        rom[603] = 12'd603;
        rom[604] = 12'd604;
        rom[605] = 12'd605;
        rom[606] = 12'd606;
        rom[607] = 12'd607;
        rom[608] = 12'd608;
        rom[609] = 12'd609;
        rom[610] = 12'd610;
        rom[611] = 12'd611;
        rom[612] = 12'd612;
        rom[613] = 12'd613;
        rom[614] = 12'd614;
        rom[615] = 12'd615;
        rom[616] = 12'd616;
        rom[617] = 12'd617;
        rom[618] = 12'd618;
        rom[619] = 12'd619;
        rom[620] = 12'd620;
        rom[621] = 12'd621;
        rom[622] = 12'd622;
        rom[623] = 12'd623;
        rom[624] = 12'd624;
        rom[625] = 12'd625;
        rom[626] = 12'd626;
        rom[627] = 12'd627;
        rom[628] = 12'd628;
        rom[629] = 12'd629;
        rom[630] = 12'd630;
        rom[631] = 12'd631;
        rom[632] = 12'd632;
        rom[633] = 12'd633;
        rom[634] = 12'd634;
        rom[635] = 12'd635;
        rom[636] = 12'd636;
        rom[637] = 12'd637;
        rom[638] = 12'd638;
        rom[639] = 12'd639;
        rom[640] = 12'd640;
        rom[641] = 12'd641;
        rom[642] = 12'd642;
        rom[643] = 12'd643;
        rom[644] = 12'd644;
        rom[645] = 12'd645;
        rom[646] = 12'd646;
        rom[647] = 12'd647;
        rom[648] = 12'd648;
        rom[649] = 12'd649;
        rom[650] = 12'd650;
        rom[651] = 12'd651;
        rom[652] = 12'd652;
        rom[653] = 12'd653;
        rom[654] = 12'd654;
        rom[655] = 12'd655;
        rom[656] = 12'd656;
        rom[657] = 12'd657;
        rom[658] = 12'd658;
        rom[659] = 12'd659;
        rom[660] = 12'd660;
        rom[661] = 12'd661;
        rom[662] = 12'd662;
        rom[663] = 12'd663;
        rom[664] = 12'd664;
        rom[665] = 12'd665;
        rom[666] = 12'd666;
        rom[667] = 12'd667;
        rom[668] = 12'd668;
        rom[669] = 12'd669;
        rom[670] = 12'd670;
        rom[671] = 12'd671;
        rom[672] = 12'd672;
        rom[673] = 12'd673;
        rom[674] = 12'd674;
        rom[675] = 12'd675;
        rom[676] = 12'd676;
        rom[677] = 12'd677;
        rom[678] = 12'd678;
        rom[679] = 12'd679;
        rom[680] = 12'd680;
        rom[681] = 12'd681;
        rom[682] = 12'd682;
        rom[683] = 12'd683;
        rom[684] = 12'd684;
        rom[685] = 12'd685;
        rom[686] = 12'd686;
        rom[687] = 12'd687;
        rom[688] = 12'd688;
        rom[689] = 12'd689;
        rom[690] = 12'd690;
        rom[691] = 12'd691;
        rom[692] = 12'd692;
        rom[693] = 12'd693;
        rom[694] = 12'd694;
        rom[695] = 12'd695;
        rom[696] = 12'd696;
        rom[697] = 12'd697;
        rom[698] = 12'd698;
        rom[699] = 12'd699;
        rom[700] = 12'd700;
        rom[701] = 12'd701;
        rom[702] = 12'd702;
        rom[703] = 12'd703;
        rom[704] = 12'd704;
        rom[705] = 12'd705;
        rom[706] = 12'd706;
        rom[707] = 12'd707;
        rom[708] = 12'd708;
        rom[709] = 12'd709;
        rom[710] = 12'd710;
        rom[711] = 12'd711;
        rom[712] = 12'd712;
        rom[713] = 12'd713;
        rom[714] = 12'd714;
        rom[715] = 12'd715;
        rom[716] = 12'd716;
        rom[717] = 12'd717;
        rom[718] = 12'd718;
        rom[719] = 12'd719;
        rom[720] = 12'd720;
        rom[721] = 12'd721;
        rom[722] = 12'd722;
        rom[723] = 12'd723;
        rom[724] = 12'd724;
        rom[725] = 12'd725;
        rom[726] = 12'd726;
        rom[727] = 12'd727;
        rom[728] = 12'd728;
        rom[729] = 12'd729;
        rom[730] = 12'd730;
        rom[731] = 12'd731;
        rom[732] = 12'd732;
        rom[733] = 12'd733;
        rom[734] = 12'd734;
        rom[735] = 12'd735;
        rom[736] = 12'd736;
        rom[737] = 12'd737;
        rom[738] = 12'd738;
        rom[739] = 12'd739;
        rom[740] = 12'd740;
        rom[741] = 12'd741;
        rom[742] = 12'd742;
        rom[743] = 12'd743;
        rom[744] = 12'd744;
        rom[745] = 12'd745;
        rom[746] = 12'd746;
        rom[747] = 12'd747;
        rom[748] = 12'd748;
        rom[749] = 12'd749;
        rom[750] = 12'd750;
        rom[751] = 12'd751;
        rom[752] = 12'd752;
        rom[753] = 12'd753;
        rom[754] = 12'd754;
        rom[755] = 12'd755;
        rom[756] = 12'd756;
        rom[757] = 12'd757;
        rom[758] = 12'd758;
        rom[759] = 12'd759;
        rom[760] = 12'd760;
        rom[761] = 12'd761;
        rom[762] = 12'd762;
        rom[763] = 12'd763;
        rom[764] = 12'd764;
        rom[765] = 12'd765;
        rom[766] = 12'd766;
        rom[767] = 12'd767;
        rom[768] = 12'd768;
        rom[769] = 12'd769;
        rom[770] = 12'd770;
        rom[771] = 12'd771;
        rom[772] = 12'd772;
        rom[773] = 12'd773;
        rom[774] = 12'd774;
        rom[775] = 12'd775;
        rom[776] = 12'd776;
        rom[777] = 12'd777;
        rom[778] = 12'd778;
        rom[779] = 12'd779;
        rom[780] = 12'd780;
        rom[781] = 12'd781;
        rom[782] = 12'd782;
        rom[783] = 12'd783;
        rom[784] = 12'd784;
        rom[785] = 12'd785;
        rom[786] = 12'd786;
        rom[787] = 12'd787;
        rom[788] = 12'd788;
        rom[789] = 12'd789;
        rom[790] = 12'd790;
        rom[791] = 12'd791;
        rom[792] = 12'd792;
        rom[793] = 12'd793;
        rom[794] = 12'd794;
        rom[795] = 12'd795;
        rom[796] = 12'd796;
        rom[797] = 12'd797;
        rom[798] = 12'd798;
        rom[799] = 12'd799;
        rom[800] = 12'd800;
        rom[801] = 12'd801;
        rom[802] = 12'd802;
        rom[803] = 12'd803;
        rom[804] = 12'd804;
        rom[805] = 12'd805;
        rom[806] = 12'd806;
        rom[807] = 12'd807;
        rom[808] = 12'd808;
        rom[809] = 12'd809;
        rom[810] = 12'd810;
        rom[811] = 12'd811;
        rom[812] = 12'd812;
        rom[813] = 12'd813;
        rom[814] = 12'd814;
        rom[815] = 12'd815;
        rom[816] = 12'd816;
        rom[817] = 12'd817;
        rom[818] = 12'd818;
        rom[819] = 12'd819;
        rom[820] = 12'd820;
        rom[821] = 12'd821;
        rom[822] = 12'd822;
        rom[823] = 12'd823;
        rom[824] = 12'd824;
        rom[825] = 12'd825;
        rom[826] = 12'd826;
        rom[827] = 12'd827;
        rom[828] = 12'd828;
        rom[829] = 12'd829;
        rom[830] = 12'd830;
        rom[831] = 12'd831;
        rom[832] = 12'd832;
        rom[833] = 12'd833;
        rom[834] = 12'd834;
        rom[835] = 12'd835;
        rom[836] = 12'd836;
        rom[837] = 12'd837;
        rom[838] = 12'd838;
        rom[839] = 12'd839;
        rom[840] = 12'd840;
        rom[841] = 12'd841;
        rom[842] = 12'd842;
        rom[843] = 12'd843;
        rom[844] = 12'd844;
        rom[845] = 12'd845;
        rom[846] = 12'd846;
        rom[847] = 12'd847;
        rom[848] = 12'd848;
        rom[849] = 12'd849;
        rom[850] = 12'd850;
        rom[851] = 12'd851;
        rom[852] = 12'd852;
        rom[853] = 12'd853;
        rom[854] = 12'd854;
        rom[855] = 12'd855;
        rom[856] = 12'd856;
        rom[857] = 12'd857;
        rom[858] = 12'd858;
        rom[859] = 12'd859;
        rom[860] = 12'd860;
        rom[861] = 12'd861;
        rom[862] = 12'd862;
        rom[863] = 12'd863;
        rom[864] = 12'd864;
        rom[865] = 12'd865;
        rom[866] = 12'd866;
        rom[867] = 12'd867;
        rom[868] = 12'd868;
        rom[869] = 12'd869;
        rom[870] = 12'd870;
        rom[871] = 12'd871;
        rom[872] = 12'd872;
        rom[873] = 12'd873;
        rom[874] = 12'd874;
        rom[875] = 12'd875;
        rom[876] = 12'd876;
        rom[877] = 12'd877;
        rom[878] = 12'd878;
        rom[879] = 12'd879;
        rom[880] = 12'd880;
        rom[881] = 12'd881;
        rom[882] = 12'd882;
        rom[883] = 12'd883;
        rom[884] = 12'd884;
        rom[885] = 12'd885;
        rom[886] = 12'd886;
        rom[887] = 12'd887;
        rom[888] = 12'd888;
        rom[889] = 12'd889;
        rom[890] = 12'd890;
        rom[891] = 12'd891;
        rom[892] = 12'd892;
        rom[893] = 12'd893;
        rom[894] = 12'd894;
        rom[895] = 12'd895;
        rom[896] = 12'd896;
        rom[897] = 12'd897;
        rom[898] = 12'd898;
        rom[899] = 12'd899;
        rom[900] = 12'd900;
        rom[901] = 12'd901;
        rom[902] = 12'd902;
        rom[903] = 12'd903;
        rom[904] = 12'd904;
        rom[905] = 12'd905;
        rom[906] = 12'd906;
        rom[907] = 12'd907;
        rom[908] = 12'd908;
        rom[909] = 12'd909;
        rom[910] = 12'd910;
        rom[911] = 12'd911;
        rom[912] = 12'd912;
        rom[913] = 12'd913;
        rom[914] = 12'd914;
        rom[915] = 12'd915;
        rom[916] = 12'd916;
        rom[917] = 12'd917;
        rom[918] = 12'd918;
        rom[919] = 12'd919;
        rom[920] = 12'd920;
        rom[921] = 12'd921;
        rom[922] = 12'd922;
        rom[923] = 12'd923;
        rom[924] = 12'd924;
        rom[925] = 12'd925;
        rom[926] = 12'd926;
        rom[927] = 12'd927;
        rom[928] = 12'd928;
        rom[929] = 12'd929;
        rom[930] = 12'd930;
        rom[931] = 12'd931;
        rom[932] = 12'd932;
        rom[933] = 12'd933;
        rom[934] = 12'd934;
        rom[935] = 12'd935;
        rom[936] = 12'd936;
        rom[937] = 12'd937;
        rom[938] = 12'd938;
        rom[939] = 12'd939;
        rom[940] = 12'd940;
        rom[941] = 12'd941;
        rom[942] = 12'd942;
        rom[943] = 12'd943;
        rom[944] = 12'd944;
        rom[945] = 12'd945;
        rom[946] = 12'd946;
        rom[947] = 12'd947;
        rom[948] = 12'd948;
        rom[949] = 12'd949;
        rom[950] = 12'd950;
        rom[951] = 12'd951;
        rom[952] = 12'd952;
        rom[953] = 12'd953;
        rom[954] = 12'd954;
        rom[955] = 12'd955;
        rom[956] = 12'd956;
        rom[957] = 12'd957;
        rom[958] = 12'd958;
        rom[959] = 12'd959;
        rom[960] = 12'd960;
        rom[961] = 12'd961;
        rom[962] = 12'd962;
        rom[963] = 12'd963;
        rom[964] = 12'd964;
        rom[965] = 12'd965;
        rom[966] = 12'd966;
        rom[967] = 12'd967;
        rom[968] = 12'd968;
        rom[969] = 12'd969;
        rom[970] = 12'd970;
        rom[971] = 12'd971;
        rom[972] = 12'd972;
        rom[973] = 12'd973;
        rom[974] = 12'd974;
        rom[975] = 12'd975;
        rom[976] = 12'd976;
        rom[977] = 12'd977;
        rom[978] = 12'd978;
        rom[979] = 12'd979;
        rom[980] = 12'd980;
        rom[981] = 12'd981;
        rom[982] = 12'd982;
        rom[983] = 12'd983;
        rom[984] = 12'd984;
        rom[985] = 12'd985;
        rom[986] = 12'd986;
        rom[987] = 12'd987;
        rom[988] = 12'd988;
        rom[989] = 12'd989;
        rom[990] = 12'd990;
        rom[991] = 12'd991;
        rom[992] = 12'd992;
        rom[993] = 12'd993;
        rom[994] = 12'd994;
        rom[995] = 12'd995;
        rom[996] = 12'd996;
        rom[997] = 12'd997;
        rom[998] = 12'd998;
        rom[999] = 12'd999;
        rom[1000] = 12'd1000;
        rom[1001] = 12'd1001;
        rom[1002] = 12'd1002;
        rom[1003] = 12'd1003;
        rom[1004] = 12'd1004;
        rom[1005] = 12'd1005;
        rom[1006] = 12'd1006;
        rom[1007] = 12'd1007;
        rom[1008] = 12'd1008;
        rom[1009] = 12'd1009;
        rom[1010] = 12'd1010;
        rom[1011] = 12'd1011;
        rom[1012] = 12'd1012;
        rom[1013] = 12'd1013;
        rom[1014] = 12'd1014;
        rom[1015] = 12'd1015;
        rom[1016] = 12'd1016;
        rom[1017] = 12'd1017;
        rom[1018] = 12'd1018;
        rom[1019] = 12'd1019;
        rom[1020] = 12'd1020;
        rom[1021] = 12'd1021;
        rom[1022] = 12'd1022;
        rom[1023] = 12'd1023;
        rom[1024] = 12'd1024;
        rom[1025] = 12'd1025;
        rom[1026] = 12'd1026;
        rom[1027] = 12'd1027;
        rom[1028] = 12'd1028;
        rom[1029] = 12'd1029;
        rom[1030] = 12'd1030;
        rom[1031] = 12'd1031;
        rom[1032] = 12'd1032;
        rom[1033] = 12'd1033;
        rom[1034] = 12'd1034;
        rom[1035] = 12'd1035;
        rom[1036] = 12'd1036;
        rom[1037] = 12'd1037;
        rom[1038] = 12'd1038;
        rom[1039] = 12'd1039;
        rom[1040] = 12'd1040;
        rom[1041] = 12'd1041;
        rom[1042] = 12'd1042;
        rom[1043] = 12'd1043;
        rom[1044] = 12'd1044;
        rom[1045] = 12'd1045;
        rom[1046] = 12'd1046;
        rom[1047] = 12'd1047;
        rom[1048] = 12'd1048;
        rom[1049] = 12'd1049;
        rom[1050] = 12'd1050;
        rom[1051] = 12'd1051;
        rom[1052] = 12'd1052;
        rom[1053] = 12'd1053;
        rom[1054] = 12'd1054;
        rom[1055] = 12'd1055;
        rom[1056] = 12'd1056;
        rom[1057] = 12'd1057;
        rom[1058] = 12'd1058;
        rom[1059] = 12'd1059;
        rom[1060] = 12'd1060;
        rom[1061] = 12'd1061;
        rom[1062] = 12'd1062;
        rom[1063] = 12'd1063;
        rom[1064] = 12'd1064;
        rom[1065] = 12'd1065;
        rom[1066] = 12'd1066;
        rom[1067] = 12'd1067;
        rom[1068] = 12'd1068;
        rom[1069] = 12'd1069;
        rom[1070] = 12'd1070;
        rom[1071] = 12'd1071;
        rom[1072] = 12'd1072;
        rom[1073] = 12'd1073;
        rom[1074] = 12'd1074;
        rom[1075] = 12'd1075;
        rom[1076] = 12'd1076;
        rom[1077] = 12'd1077;
        rom[1078] = 12'd1078;
        rom[1079] = 12'd1079;
        rom[1080] = 12'd1080;
        rom[1081] = 12'd1081;
        rom[1082] = 12'd1082;
        rom[1083] = 12'd1083;
        rom[1084] = 12'd1084;
        rom[1085] = 12'd1085;
        rom[1086] = 12'd1086;
        rom[1087] = 12'd1087;
        rom[1088] = 12'd1088;
        rom[1089] = 12'd1089;
        rom[1090] = 12'd1090;
        rom[1091] = 12'd1091;
        rom[1092] = 12'd1092;
        rom[1093] = 12'd1093;
        rom[1094] = 12'd1094;
        rom[1095] = 12'd1095;
        rom[1096] = 12'd1096;
        rom[1097] = 12'd1097;
        rom[1098] = 12'd1098;
        rom[1099] = 12'd1099;
        rom[1100] = 12'd1100;
        rom[1101] = 12'd1101;
        rom[1102] = 12'd1102;
        rom[1103] = 12'd1103;
        rom[1104] = 12'd1104;
        rom[1105] = 12'd1105;
        rom[1106] = 12'd1106;
        rom[1107] = 12'd1107;
        rom[1108] = 12'd1108;
        rom[1109] = 12'd1109;
        rom[1110] = 12'd1110;
        rom[1111] = 12'd1111;
        rom[1112] = 12'd1112;
        rom[1113] = 12'd1113;
        rom[1114] = 12'd1114;
        rom[1115] = 12'd1115;
        rom[1116] = 12'd1116;
        rom[1117] = 12'd1117;
        rom[1118] = 12'd1118;
        rom[1119] = 12'd1119;
        rom[1120] = 12'd1120;
        rom[1121] = 12'd1121;
        rom[1122] = 12'd1122;
        rom[1123] = 12'd1123;
        rom[1124] = 12'd1124;
        rom[1125] = 12'd1125;
        rom[1126] = 12'd1126;
        rom[1127] = 12'd1127;
        rom[1128] = 12'd1128;
        rom[1129] = 12'd1129;
        rom[1130] = 12'd1130;
        rom[1131] = 12'd1131;
        rom[1132] = 12'd1132;
        rom[1133] = 12'd1133;
        rom[1134] = 12'd1134;
        rom[1135] = 12'd1135;
        rom[1136] = 12'd1136;
        rom[1137] = 12'd1137;
        rom[1138] = 12'd1138;
        rom[1139] = 12'd1139;
        rom[1140] = 12'd1140;
        rom[1141] = 12'd1141;
        rom[1142] = 12'd1142;
        rom[1143] = 12'd1143;
        rom[1144] = 12'd1144;
        rom[1145] = 12'd1145;
        rom[1146] = 12'd1146;
        rom[1147] = 12'd1147;
        rom[1148] = 12'd1148;
        rom[1149] = 12'd1149;
        rom[1150] = 12'd1150;
        rom[1151] = 12'd1151;
        rom[1152] = 12'd1152;
        rom[1153] = 12'd1153;
        rom[1154] = 12'd1154;
        rom[1155] = 12'd1155;
        rom[1156] = 12'd1156;
        rom[1157] = 12'd1157;
        rom[1158] = 12'd1158;
        rom[1159] = 12'd1159;
        rom[1160] = 12'd1160;
        rom[1161] = 12'd1161;
        rom[1162] = 12'd1162;
        rom[1163] = 12'd1163;
        rom[1164] = 12'd1164;
        rom[1165] = 12'd1165;
        rom[1166] = 12'd1166;
        rom[1167] = 12'd1167;
        rom[1168] = 12'd1168;
        rom[1169] = 12'd1169;
        rom[1170] = 12'd1170;
        rom[1171] = 12'd1171;
        rom[1172] = 12'd1172;
        rom[1173] = 12'd1173;
        rom[1174] = 12'd1174;
        rom[1175] = 12'd1175;
        rom[1176] = 12'd1176;
        rom[1177] = 12'd1177;
        rom[1178] = 12'd1178;
        rom[1179] = 12'd1179;
        rom[1180] = 12'd1180;
        rom[1181] = 12'd1181;
        rom[1182] = 12'd1182;
        rom[1183] = 12'd1183;
        rom[1184] = 12'd1184;
        rom[1185] = 12'd1185;
        rom[1186] = 12'd1186;
        rom[1187] = 12'd1187;
        rom[1188] = 12'd1188;
        rom[1189] = 12'd1189;
        rom[1190] = 12'd1190;
        rom[1191] = 12'd1191;
        rom[1192] = 12'd1192;
        rom[1193] = 12'd1193;
        rom[1194] = 12'd1194;
        rom[1195] = 12'd1195;
        rom[1196] = 12'd1196;
        rom[1197] = 12'd1197;
        rom[1198] = 12'd1198;
        rom[1199] = 12'd1199;
        rom[1200] = 12'd1200;
        rom[1201] = 12'd1201;
        rom[1202] = 12'd1202;
        rom[1203] = 12'd1203;
        rom[1204] = 12'd1204;
        rom[1205] = 12'd1205;
        rom[1206] = 12'd1206;
        rom[1207] = 12'd1207;
        rom[1208] = 12'd1208;
        rom[1209] = 12'd1209;
        rom[1210] = 12'd1210;
        rom[1211] = 12'd1211;
        rom[1212] = 12'd1212;
        rom[1213] = 12'd1213;
        rom[1214] = 12'd1214;
        rom[1215] = 12'd1215;
        rom[1216] = 12'd1216;
        rom[1217] = 12'd1217;
        rom[1218] = 12'd1218;
        rom[1219] = 12'd1219;
        rom[1220] = 12'd1220;
        rom[1221] = 12'd1221;
        rom[1222] = 12'd1222;
        rom[1223] = 12'd1223;
        rom[1224] = 12'd1224;
        rom[1225] = 12'd1225;
        rom[1226] = 12'd1226;
        rom[1227] = 12'd1227;
        rom[1228] = 12'd1228;
        rom[1229] = 12'd1229;
        rom[1230] = 12'd1230;
        rom[1231] = 12'd1231;
        rom[1232] = 12'd1232;
        rom[1233] = 12'd1233;
        rom[1234] = 12'd1234;
        rom[1235] = 12'd1235;
        rom[1236] = 12'd1236;
        rom[1237] = 12'd1237;
        rom[1238] = 12'd1238;
        rom[1239] = 12'd1239;
        rom[1240] = 12'd1240;
        rom[1241] = 12'd1241;
        rom[1242] = 12'd1242;
        rom[1243] = 12'd1243;
        rom[1244] = 12'd1244;
        rom[1245] = 12'd1245;
        rom[1246] = 12'd1246;
        rom[1247] = 12'd1247;
        rom[1248] = 12'd1248;
        rom[1249] = 12'd1249;
        rom[1250] = 12'd1250;
        rom[1251] = 12'd1251;
        rom[1252] = 12'd1252;
        rom[1253] = 12'd1253;
        rom[1254] = 12'd1254;
        rom[1255] = 12'd1255;
        rom[1256] = 12'd1256;
        rom[1257] = 12'd1257;
        rom[1258] = 12'd1258;
        rom[1259] = 12'd1259;
        rom[1260] = 12'd1260;
        rom[1261] = 12'd1261;
        rom[1262] = 12'd1262;
        rom[1263] = 12'd1263;
        rom[1264] = 12'd1264;
        rom[1265] = 12'd1265;
        rom[1266] = 12'd1266;
        rom[1267] = 12'd1267;
        rom[1268] = 12'd1268;
        rom[1269] = 12'd1269;
        rom[1270] = 12'd1270;
        rom[1271] = 12'd1271;
        rom[1272] = 12'd1272;
        rom[1273] = 12'd1273;
        rom[1274] = 12'd1274;
        rom[1275] = 12'd1275;
        rom[1276] = 12'd1276;
        rom[1277] = 12'd1277;
        rom[1278] = 12'd1278;
        rom[1279] = 12'd1279;
        rom[1280] = 12'd1280;
        rom[1281] = 12'd1281;
        rom[1282] = 12'd1282;
        rom[1283] = 12'd1283;
        rom[1284] = 12'd1284;
        rom[1285] = 12'd1285;
        rom[1286] = 12'd1286;
        rom[1287] = 12'd1287;
        rom[1288] = 12'd1288;
        rom[1289] = 12'd1289;
        rom[1290] = 12'd1290;
        rom[1291] = 12'd1291;
        rom[1292] = 12'd1292;
        rom[1293] = 12'd1293;
        rom[1294] = 12'd1294;
        rom[1295] = 12'd1295;
        rom[1296] = 12'd1296;
        rom[1297] = 12'd1297;
        rom[1298] = 12'd1298;
        rom[1299] = 12'd1299;
        rom[1300] = 12'd1300;
        rom[1301] = 12'd1301;
        rom[1302] = 12'd1302;
        rom[1303] = 12'd1303;
        rom[1304] = 12'd1304;
        rom[1305] = 12'd1305;
        rom[1306] = 12'd1306;
        rom[1307] = 12'd1307;
        rom[1308] = 12'd1308;
        rom[1309] = 12'd1309;
        rom[1310] = 12'd1310;
        rom[1311] = 12'd1311;
        rom[1312] = 12'd1312;
        rom[1313] = 12'd1313;
        rom[1314] = 12'd1314;
        rom[1315] = 12'd1315;
        rom[1316] = 12'd1316;
        rom[1317] = 12'd1317;
        rom[1318] = 12'd1318;
        rom[1319] = 12'd1319;
        rom[1320] = 12'd1320;
        rom[1321] = 12'd1321;
        rom[1322] = 12'd1322;
        rom[1323] = 12'd1323;
        rom[1324] = 12'd1324;
        rom[1325] = 12'd1325;
        rom[1326] = 12'd1326;
        rom[1327] = 12'd1327;
        rom[1328] = 12'd1328;
        rom[1329] = 12'd1329;
        rom[1330] = 12'd1330;
        rom[1331] = 12'd1331;
        rom[1332] = 12'd1332;
        rom[1333] = 12'd1333;
        rom[1334] = 12'd1334;
        rom[1335] = 12'd1335;
        rom[1336] = 12'd1336;
        rom[1337] = 12'd1337;
        rom[1338] = 12'd1338;
        rom[1339] = 12'd1339;
        rom[1340] = 12'd1340;
        rom[1341] = 12'd1341;
        rom[1342] = 12'd1342;
        rom[1343] = 12'd1343;
        rom[1344] = 12'd1344;
        rom[1345] = 12'd1345;
        rom[1346] = 12'd1346;
        rom[1347] = 12'd1347;
        rom[1348] = 12'd1348;
        rom[1349] = 12'd1349;
        rom[1350] = 12'd1350;
        rom[1351] = 12'd1351;
        rom[1352] = 12'd1352;
        rom[1353] = 12'd1353;
        rom[1354] = 12'd1354;
        rom[1355] = 12'd1355;
        rom[1356] = 12'd1356;
        rom[1357] = 12'd1357;
        rom[1358] = 12'd1358;
        rom[1359] = 12'd1359;
        rom[1360] = 12'd1360;
        rom[1361] = 12'd1361;
        rom[1362] = 12'd1362;
        rom[1363] = 12'd1363;
        rom[1364] = 12'd1364;
        rom[1365] = 12'd1365;
        rom[1366] = 12'd1366;
        rom[1367] = 12'd1367;
        rom[1368] = 12'd1368;
        rom[1369] = 12'd1369;
        rom[1370] = 12'd1370;
        rom[1371] = 12'd1371;
        rom[1372] = 12'd1372;
        rom[1373] = 12'd1373;
        rom[1374] = 12'd1374;
        rom[1375] = 12'd1375;
        rom[1376] = 12'd1376;
        rom[1377] = 12'd1377;
        rom[1378] = 12'd1378;
        rom[1379] = 12'd1379;
        rom[1380] = 12'd1380;
        rom[1381] = 12'd1381;
        rom[1382] = 12'd1382;
        rom[1383] = 12'd1383;
        rom[1384] = 12'd1384;
        rom[1385] = 12'd1385;
        rom[1386] = 12'd1386;
        rom[1387] = 12'd1387;
        rom[1388] = 12'd1388;
        rom[1389] = 12'd1389;
        rom[1390] = 12'd1390;
        rom[1391] = 12'd1391;
        rom[1392] = 12'd1392;
        rom[1393] = 12'd1393;
        rom[1394] = 12'd1394;
        rom[1395] = 12'd1395;
        rom[1396] = 12'd1396;
        rom[1397] = 12'd1397;
        rom[1398] = 12'd1398;
        rom[1399] = 12'd1399;
        rom[1400] = 12'd1400;
        rom[1401] = 12'd1401;
        rom[1402] = 12'd1402;
        rom[1403] = 12'd1403;
        rom[1404] = 12'd1404;
        rom[1405] = 12'd1405;
        rom[1406] = 12'd1406;
        rom[1407] = 12'd1407;
        rom[1408] = 12'd1408;
        rom[1409] = 12'd1409;
        rom[1410] = 12'd1410;
        rom[1411] = 12'd1411;
        rom[1412] = 12'd1412;
        rom[1413] = 12'd1413;
        rom[1414] = 12'd1414;
        rom[1415] = 12'd1415;
        rom[1416] = 12'd1416;
        rom[1417] = 12'd1417;
        rom[1418] = 12'd1418;
        rom[1419] = 12'd1419;
        rom[1420] = 12'd1420;
        rom[1421] = 12'd1421;
        rom[1422] = 12'd1422;
        rom[1423] = 12'd1423;
        rom[1424] = 12'd1424;
        rom[1425] = 12'd1425;
        rom[1426] = 12'd1426;
        rom[1427] = 12'd1427;
        rom[1428] = 12'd1428;
        rom[1429] = 12'd1429;
        rom[1430] = 12'd1430;
        rom[1431] = 12'd1431;
        rom[1432] = 12'd1432;
        rom[1433] = 12'd1433;
        rom[1434] = 12'd1434;
        rom[1435] = 12'd1435;
        rom[1436] = 12'd1436;
        rom[1437] = 12'd1437;
        rom[1438] = 12'd1438;
        rom[1439] = 12'd1439;
        rom[1440] = 12'd1440;
        rom[1441] = 12'd1441;
        rom[1442] = 12'd1442;
        rom[1443] = 12'd1443;
        rom[1444] = 12'd1444;
        rom[1445] = 12'd1445;
        rom[1446] = 12'd1446;
        rom[1447] = 12'd1447;
        rom[1448] = 12'd1448;
        rom[1449] = 12'd1449;
        rom[1450] = 12'd1450;
        rom[1451] = 12'd1451;
        rom[1452] = 12'd1452;
        rom[1453] = 12'd1453;
        rom[1454] = 12'd1454;
        rom[1455] = 12'd1455;
        rom[1456] = 12'd1456;
        rom[1457] = 12'd1457;
        rom[1458] = 12'd1458;
        rom[1459] = 12'd1459;
        rom[1460] = 12'd1460;
        rom[1461] = 12'd1461;
        rom[1462] = 12'd1462;
        rom[1463] = 12'd1463;
        rom[1464] = 12'd1464;
        rom[1465] = 12'd1465;
        rom[1466] = 12'd1466;
        rom[1467] = 12'd1467;
        rom[1468] = 12'd1468;
        rom[1469] = 12'd1469;
        rom[1470] = 12'd1470;
        rom[1471] = 12'd1471;
        rom[1472] = 12'd1472;
        rom[1473] = 12'd1473;
        rom[1474] = 12'd1474;
        rom[1475] = 12'd1475;
        rom[1476] = 12'd1476;
        rom[1477] = 12'd1477;
        rom[1478] = 12'd1478;
        rom[1479] = 12'd1479;
        rom[1480] = 12'd1480;
        rom[1481] = 12'd1481;
        rom[1482] = 12'd1482;
        rom[1483] = 12'd1483;
        rom[1484] = 12'd1484;
        rom[1485] = 12'd1485;
        rom[1486] = 12'd1486;
        rom[1487] = 12'd1487;
        rom[1488] = 12'd1488;
        rom[1489] = 12'd1489;
        rom[1490] = 12'd1490;
        rom[1491] = 12'd1491;
        rom[1492] = 12'd1492;
        rom[1493] = 12'd1493;
        rom[1494] = 12'd1494;
        rom[1495] = 12'd1495;
        rom[1496] = 12'd1496;
        rom[1497] = 12'd1497;
        rom[1498] = 12'd1498;
        rom[1499] = 12'd1499;
        rom[1500] = 12'd1500;
        rom[1501] = 12'd1501;
        rom[1502] = 12'd1502;
        rom[1503] = 12'd1503;
        rom[1504] = 12'd1504;
        rom[1505] = 12'd1505;
        rom[1506] = 12'd1506;
        rom[1507] = 12'd1507;
        rom[1508] = 12'd1508;
        rom[1509] = 12'd1509;
        rom[1510] = 12'd1510;
        rom[1511] = 12'd1511;
        rom[1512] = 12'd1512;
        rom[1513] = 12'd1513;
        rom[1514] = 12'd1514;
        rom[1515] = 12'd1515;
        rom[1516] = 12'd1516;
        rom[1517] = 12'd1517;
        rom[1518] = 12'd1518;
        rom[1519] = 12'd1519;
        rom[1520] = 12'd1520;
        rom[1521] = 12'd1521;
        rom[1522] = 12'd1522;
        rom[1523] = 12'd1523;
        rom[1524] = 12'd1524;
        rom[1525] = 12'd1525;
        rom[1526] = 12'd1526;
        rom[1527] = 12'd1527;
        rom[1528] = 12'd1528;
        rom[1529] = 12'd1529;
        rom[1530] = 12'd1530;
        rom[1531] = 12'd1531;
        rom[1532] = 12'd1532;
        rom[1533] = 12'd1533;
        rom[1534] = 12'd1534;
        rom[1535] = 12'd1535;
        rom[1536] = 12'd1536;
        rom[1537] = 12'd1537;
        rom[1538] = 12'd1538;
        rom[1539] = 12'd1539;
        rom[1540] = 12'd1540;
        rom[1541] = 12'd1541;
        rom[1542] = 12'd1542;
        rom[1543] = 12'd1543;
        rom[1544] = 12'd1544;
        rom[1545] = 12'd1545;
        rom[1546] = 12'd1546;
        rom[1547] = 12'd1547;
        rom[1548] = 12'd1548;
        rom[1549] = 12'd1549;
        rom[1550] = 12'd1550;
        rom[1551] = 12'd1551;
        rom[1552] = 12'd1552;
        rom[1553] = 12'd1553;
        rom[1554] = 12'd1554;
        rom[1555] = 12'd1555;
        rom[1556] = 12'd1556;
        rom[1557] = 12'd1557;
        rom[1558] = 12'd1558;
        rom[1559] = 12'd1559;
        rom[1560] = 12'd1560;
        rom[1561] = 12'd1561;
        rom[1562] = 12'd1562;
        rom[1563] = 12'd1563;
        rom[1564] = 12'd1564;
        rom[1565] = 12'd1565;
        rom[1566] = 12'd1566;
        rom[1567] = 12'd1567;
        rom[1568] = 12'd1568;
        rom[1569] = 12'd1569;
        rom[1570] = 12'd1570;
        rom[1571] = 12'd1571;
        rom[1572] = 12'd1572;
        rom[1573] = 12'd1573;
        rom[1574] = 12'd1574;
        rom[1575] = 12'd1575;
        rom[1576] = 12'd1576;
        rom[1577] = 12'd1577;
        rom[1578] = 12'd1578;
        rom[1579] = 12'd1579;
        rom[1580] = 12'd1580;
        rom[1581] = 12'd1581;
        rom[1582] = 12'd1582;
        rom[1583] = 12'd1583;
        rom[1584] = 12'd1584;
        rom[1585] = 12'd1585;
        rom[1586] = 12'd1586;
        rom[1587] = 12'd1587;
        rom[1588] = 12'd1588;
        rom[1589] = 12'd1589;
        rom[1590] = 12'd1590;
        rom[1591] = 12'd1591;
        rom[1592] = 12'd1592;
        rom[1593] = 12'd1593;
        rom[1594] = 12'd1594;
        rom[1595] = 12'd1595;
        rom[1596] = 12'd1596;
        rom[1597] = 12'd1597;
        rom[1598] = 12'd1598;
        rom[1599] = 12'd1599;
        rom[1600] = 12'd1600;
        rom[1601] = 12'd1601;
        rom[1602] = 12'd1602;
        rom[1603] = 12'd1603;
        rom[1604] = 12'd1604;
        rom[1605] = 12'd1605;
        rom[1606] = 12'd1606;
        rom[1607] = 12'd1607;
        rom[1608] = 12'd1608;
        rom[1609] = 12'd1609;
        rom[1610] = 12'd1610;
        rom[1611] = 12'd1611;
        rom[1612] = 12'd1612;
        rom[1613] = 12'd1613;
        rom[1614] = 12'd1614;
        rom[1615] = 12'd1615;
        rom[1616] = 12'd1616;
        rom[1617] = 12'd1617;
        rom[1618] = 12'd1618;
        rom[1619] = 12'd1619;
        rom[1620] = 12'd1620;
        rom[1621] = 12'd1621;
        rom[1622] = 12'd1622;
        rom[1623] = 12'd1623;
        rom[1624] = 12'd1624;
        rom[1625] = 12'd1625;
        rom[1626] = 12'd1626;
        rom[1627] = 12'd1627;
        rom[1628] = 12'd1628;
        rom[1629] = 12'd1629;
        rom[1630] = 12'd1630;
        rom[1631] = 12'd1631;
        rom[1632] = 12'd1632;
        rom[1633] = 12'd1633;
        rom[1634] = 12'd1634;
        rom[1635] = 12'd1635;
        rom[1636] = 12'd1636;
        rom[1637] = 12'd1637;
        rom[1638] = 12'd1638;
        rom[1639] = 12'd1639;
        rom[1640] = 12'd1640;
        rom[1641] = 12'd1641;
        rom[1642] = 12'd1642;
        rom[1643] = 12'd1643;
        rom[1644] = 12'd1644;
        rom[1645] = 12'd1645;
        rom[1646] = 12'd1646;
        rom[1647] = 12'd1647;
        rom[1648] = 12'd1648;
        rom[1649] = 12'd1649;
        rom[1650] = 12'd1650;
        rom[1651] = 12'd1651;
        rom[1652] = 12'd1652;
        rom[1653] = 12'd1653;
        rom[1654] = 12'd1654;
        rom[1655] = 12'd1655;
        rom[1656] = 12'd1656;
        rom[1657] = 12'd1657;
        rom[1658] = 12'd1658;
        rom[1659] = 12'd1659;
        rom[1660] = 12'd1660;
        rom[1661] = 12'd1661;
        rom[1662] = 12'd1662;
        rom[1663] = 12'd1663;
        rom[1664] = 12'd1664;
        rom[1665] = 12'd1665;
        rom[1666] = 12'd1666;
        rom[1667] = 12'd1667;
        rom[1668] = 12'd1668;
        rom[1669] = 12'd1669;
        rom[1670] = 12'd1670;
        rom[1671] = 12'd1671;
        rom[1672] = 12'd1672;
        rom[1673] = 12'd1673;
        rom[1674] = 12'd1674;
        rom[1675] = 12'd1675;
        rom[1676] = 12'd1676;
        rom[1677] = 12'd1677;
        rom[1678] = 12'd1678;
        rom[1679] = 12'd1679;
        rom[1680] = 12'd1680;
        rom[1681] = 12'd1681;
        rom[1682] = 12'd1682;
        rom[1683] = 12'd1683;
        rom[1684] = 12'd1684;
        rom[1685] = 12'd1685;
        rom[1686] = 12'd1686;
        rom[1687] = 12'd1687;
        rom[1688] = 12'd1688;
        rom[1689] = 12'd1689;
        rom[1690] = 12'd1690;
        rom[1691] = 12'd1691;
        rom[1692] = 12'd1692;
        rom[1693] = 12'd1693;
        rom[1694] = 12'd1694;
        rom[1695] = 12'd1695;
        rom[1696] = 12'd1696;
        rom[1697] = 12'd1697;
        rom[1698] = 12'd1698;
        rom[1699] = 12'd1699;
        rom[1700] = 12'd1700;
        rom[1701] = 12'd1701;
        rom[1702] = 12'd1702;
        rom[1703] = 12'd1703;
        rom[1704] = 12'd1704;
        rom[1705] = 12'd1705;
        rom[1706] = 12'd1706;
        rom[1707] = 12'd1707;
        rom[1708] = 12'd1708;
        rom[1709] = 12'd1709;
        rom[1710] = 12'd1710;
        rom[1711] = 12'd1711;
        rom[1712] = 12'd1712;
        rom[1713] = 12'd1713;
        rom[1714] = 12'd1714;
        rom[1715] = 12'd1715;
        rom[1716] = 12'd1716;
        rom[1717] = 12'd1717;
        rom[1718] = 12'd1718;
        rom[1719] = 12'd1719;
        rom[1720] = 12'd1720;
        rom[1721] = 12'd1721;
        rom[1722] = 12'd1722;
        rom[1723] = 12'd1723;
        rom[1724] = 12'd1724;
        rom[1725] = 12'd1725;
        rom[1726] = 12'd1726;
        rom[1727] = 12'd1727;
        rom[1728] = 12'd1728;
        rom[1729] = 12'd1729;
        rom[1730] = 12'd1730;
        rom[1731] = 12'd1731;
        rom[1732] = 12'd1732;
        rom[1733] = 12'd1733;
        rom[1734] = 12'd1734;
        rom[1735] = 12'd1735;
        rom[1736] = 12'd1736;
        rom[1737] = 12'd1737;
        rom[1738] = 12'd1738;
        rom[1739] = 12'd1739;
        rom[1740] = 12'd1740;
        rom[1741] = 12'd1741;
        rom[1742] = 12'd1742;
        rom[1743] = 12'd1743;
        rom[1744] = 12'd1744;
        rom[1745] = 12'd1745;
        rom[1746] = 12'd1746;
        rom[1747] = 12'd1747;
        rom[1748] = 12'd1748;
        rom[1749] = 12'd1749;
        rom[1750] = 12'd1750;
        rom[1751] = 12'd1751;
        rom[1752] = 12'd1752;
        rom[1753] = 12'd1753;
        rom[1754] = 12'd1754;
        rom[1755] = 12'd1755;
        rom[1756] = 12'd1756;
        rom[1757] = 12'd1757;
        rom[1758] = 12'd1758;
        rom[1759] = 12'd1759;
        rom[1760] = 12'd1760;
        rom[1761] = 12'd1761;
        rom[1762] = 12'd1762;
        rom[1763] = 12'd1763;
        rom[1764] = 12'd1764;
        rom[1765] = 12'd1765;
        rom[1766] = 12'd1766;
        rom[1767] = 12'd1767;
        rom[1768] = 12'd1768;
        rom[1769] = 12'd1769;
        rom[1770] = 12'd1770;
        rom[1771] = 12'd1771;
        rom[1772] = 12'd1772;
        rom[1773] = 12'd1773;
        rom[1774] = 12'd1774;
        rom[1775] = 12'd1775;
        rom[1776] = 12'd1776;
        rom[1777] = 12'd1777;
        rom[1778] = 12'd1778;
        rom[1779] = 12'd1779;
        rom[1780] = 12'd1780;
        rom[1781] = 12'd1781;
        rom[1782] = 12'd1782;
        rom[1783] = 12'd1783;
        rom[1784] = 12'd1784;
        rom[1785] = 12'd1785;
        rom[1786] = 12'd1786;
        rom[1787] = 12'd1787;
        rom[1788] = 12'd1788;
        rom[1789] = 12'd1789;
        rom[1790] = 12'd1790;
        rom[1791] = 12'd1791;
        rom[1792] = 12'd1792;
        rom[1793] = 12'd1793;
        rom[1794] = 12'd1794;
        rom[1795] = 12'd1795;
        rom[1796] = 12'd1796;
        rom[1797] = 12'd1797;
        rom[1798] = 12'd1798;
        rom[1799] = 12'd1799;
        rom[1800] = 12'd1800;
        rom[1801] = 12'd1801;
        rom[1802] = 12'd1802;
        rom[1803] = 12'd1803;
        rom[1804] = 12'd1804;
        rom[1805] = 12'd1805;
        rom[1806] = 12'd1806;
        rom[1807] = 12'd1807;
        rom[1808] = 12'd1808;
        rom[1809] = 12'd1809;
        rom[1810] = 12'd1810;
        rom[1811] = 12'd1811;
        rom[1812] = 12'd1812;
        rom[1813] = 12'd1813;
        rom[1814] = 12'd1814;
        rom[1815] = 12'd1815;
        rom[1816] = 12'd1816;
        rom[1817] = 12'd1817;
        rom[1818] = 12'd1818;
        rom[1819] = 12'd1819;
        rom[1820] = 12'd1820;
        rom[1821] = 12'd1821;
        rom[1822] = 12'd1822;
        rom[1823] = 12'd1823;
        rom[1824] = 12'd1824;
        rom[1825] = 12'd1825;
        rom[1826] = 12'd1826;
        rom[1827] = 12'd1827;
        rom[1828] = 12'd1828;
        rom[1829] = 12'd1829;
        rom[1830] = 12'd1830;
        rom[1831] = 12'd1831;
        rom[1832] = 12'd1832;
        rom[1833] = 12'd1833;
        rom[1834] = 12'd1834;
        rom[1835] = 12'd1835;
        rom[1836] = 12'd1836;
        rom[1837] = 12'd1837;
        rom[1838] = 12'd1838;
        rom[1839] = 12'd1839;
        rom[1840] = 12'd1840;
        rom[1841] = 12'd1841;
        rom[1842] = 12'd1842;
        rom[1843] = 12'd1843;
        rom[1844] = 12'd1844;
        rom[1845] = 12'd1845;
        rom[1846] = 12'd1846;
        rom[1847] = 12'd1847;
        rom[1848] = 12'd1848;
        rom[1849] = 12'd1849;
        rom[1850] = 12'd1850;
        rom[1851] = 12'd1851;
        rom[1852] = 12'd1852;
        rom[1853] = 12'd1853;
        rom[1854] = 12'd1854;
        rom[1855] = 12'd1855;
        rom[1856] = 12'd1856;
        rom[1857] = 12'd1857;
        rom[1858] = 12'd1858;
        rom[1859] = 12'd1859;
        rom[1860] = 12'd1860;
        rom[1861] = 12'd1861;
        rom[1862] = 12'd1862;
        rom[1863] = 12'd1863;
        rom[1864] = 12'd1864;
        rom[1865] = 12'd1865;
        rom[1866] = 12'd1866;
        rom[1867] = 12'd1867;
        rom[1868] = 12'd1868;
        rom[1869] = 12'd1869;
        rom[1870] = 12'd1870;
        rom[1871] = 12'd1871;
        rom[1872] = 12'd1872;
        rom[1873] = 12'd1873;
        rom[1874] = 12'd1874;
        rom[1875] = 12'd1875;
        rom[1876] = 12'd1876;
        rom[1877] = 12'd1877;
        rom[1878] = 12'd1878;
        rom[1879] = 12'd1879;
        rom[1880] = 12'd1880;
        rom[1881] = 12'd1881;
        rom[1882] = 12'd1882;
        rom[1883] = 12'd1883;
        rom[1884] = 12'd1884;
        rom[1885] = 12'd1885;
        rom[1886] = 12'd1886;
        rom[1887] = 12'd1887;
        rom[1888] = 12'd1888;
        rom[1889] = 12'd1889;
        rom[1890] = 12'd1890;
        rom[1891] = 12'd1891;
        rom[1892] = 12'd1892;
        rom[1893] = 12'd1893;
        rom[1894] = 12'd1894;
        rom[1895] = 12'd1895;
        rom[1896] = 12'd1896;
        rom[1897] = 12'd1897;
        rom[1898] = 12'd1898;
        rom[1899] = 12'd1899;
        rom[1900] = 12'd1900;
        rom[1901] = 12'd1901;
        rom[1902] = 12'd1902;
        rom[1903] = 12'd1903;
        rom[1904] = 12'd1904;
        rom[1905] = 12'd1905;
        rom[1906] = 12'd1906;
        rom[1907] = 12'd1907;
        rom[1908] = 12'd1908;
        rom[1909] = 12'd1909;
        rom[1910] = 12'd1910;
        rom[1911] = 12'd1911;
        rom[1912] = 12'd1912;
        rom[1913] = 12'd1913;
        rom[1914] = 12'd1914;
        rom[1915] = 12'd1915;
        rom[1916] = 12'd1916;
        rom[1917] = 12'd1917;
        rom[1918] = 12'd1918;
        rom[1919] = 12'd1919;
        rom[1920] = 12'd1920;
        rom[1921] = 12'd1921;
        rom[1922] = 12'd1922;
        rom[1923] = 12'd1923;
        rom[1924] = 12'd1924;
        rom[1925] = 12'd1925;
        rom[1926] = 12'd1926;
        rom[1927] = 12'd1927;
        rom[1928] = 12'd1928;
        rom[1929] = 12'd1929;
        rom[1930] = 12'd1930;
        rom[1931] = 12'd1931;
        rom[1932] = 12'd1932;
        rom[1933] = 12'd1933;
        rom[1934] = 12'd1934;
        rom[1935] = 12'd1935;
        rom[1936] = 12'd1936;
        rom[1937] = 12'd1937;
        rom[1938] = 12'd1938;
        rom[1939] = 12'd1939;
        rom[1940] = 12'd1940;
        rom[1941] = 12'd1941;
        rom[1942] = 12'd1942;
        rom[1943] = 12'd1943;
        rom[1944] = 12'd1944;
        rom[1945] = 12'd1945;
        rom[1946] = 12'd1946;
        rom[1947] = 12'd1947;
        rom[1948] = 12'd1948;
        rom[1949] = 12'd1949;
        rom[1950] = 12'd1950;
        rom[1951] = 12'd1951;
        rom[1952] = 12'd1952;
        rom[1953] = 12'd1953;
        rom[1954] = 12'd1954;
        rom[1955] = 12'd1955;
        rom[1956] = 12'd1956;
        rom[1957] = 12'd1957;
        rom[1958] = 12'd1958;
        rom[1959] = 12'd1959;
        rom[1960] = 12'd1960;
        rom[1961] = 12'd1961;
        rom[1962] = 12'd1962;
        rom[1963] = 12'd1963;
        rom[1964] = 12'd1964;
        rom[1965] = 12'd1965;
        rom[1966] = 12'd1966;
        rom[1967] = 12'd1967;
        rom[1968] = 12'd1968;
        rom[1969] = 12'd1969;
        rom[1970] = 12'd1970;
        rom[1971] = 12'd1971;
        rom[1972] = 12'd1972;
        rom[1973] = 12'd1973;
        rom[1974] = 12'd1974;
        rom[1975] = 12'd1975;
        rom[1976] = 12'd1976;
        rom[1977] = 12'd1977;
        rom[1978] = 12'd1978;
        rom[1979] = 12'd1979;
        rom[1980] = 12'd1980;
        rom[1981] = 12'd1981;
        rom[1982] = 12'd1982;
        rom[1983] = 12'd1983;
        rom[1984] = 12'd1984;
        rom[1985] = 12'd1985;
        rom[1986] = 12'd1986;
        rom[1987] = 12'd1987;
        rom[1988] = 12'd1988;
        rom[1989] = 12'd1989;
        rom[1990] = 12'd1990;
        rom[1991] = 12'd1991;
        rom[1992] = 12'd1992;
        rom[1993] = 12'd1993;
        rom[1994] = 12'd1994;
        rom[1995] = 12'd1995;
        rom[1996] = 12'd1996;
        rom[1997] = 12'd1997;
        rom[1998] = 12'd1998;
        rom[1999] = 12'd1999;
        rom[2000] = 12'd2000;
        rom[2001] = 12'd2001;
        rom[2002] = 12'd2002;
        rom[2003] = 12'd2003;
        rom[2004] = 12'd2004;
        rom[2005] = 12'd2005;
        rom[2006] = 12'd2006;
        rom[2007] = 12'd2007;
        rom[2008] = 12'd2008;
        rom[2009] = 12'd2009;
        rom[2010] = 12'd2010;
        rom[2011] = 12'd2011;
        rom[2012] = 12'd2012;
        rom[2013] = 12'd2013;
        rom[2014] = 12'd2014;
        rom[2015] = 12'd2015;
        rom[2016] = 12'd2016;
        rom[2017] = 12'd2017;
        rom[2018] = 12'd2018;
        rom[2019] = 12'd2019;
        rom[2020] = 12'd2020;
        rom[2021] = 12'd2021;
        rom[2022] = 12'd2022;
        rom[2023] = 12'd2023;
        rom[2024] = 12'd2024;
        rom[2025] = 12'd2025;
        rom[2026] = 12'd2026;
        rom[2027] = 12'd2027;
        rom[2028] = 12'd2028;
        rom[2029] = 12'd2029;
        rom[2030] = 12'd2030;
        rom[2031] = 12'd2031;
        rom[2032] = 12'd2032;
        rom[2033] = 12'd2033;
        rom[2034] = 12'd2034;
        rom[2035] = 12'd2035;
        rom[2036] = 12'd2036;
        rom[2037] = 12'd2037;
        rom[2038] = 12'd2038;
        rom[2039] = 12'd2039;
        rom[2040] = 12'd2040;
        rom[2041] = 12'd2041;
        rom[2042] = 12'd2042;
        rom[2043] = 12'd2043;
        rom[2044] = 12'd2044;
        rom[2045] = 12'd2045;
        rom[2046] = 12'd2046;
        rom[2047] = 12'd2047;
        rom[2048] = 12'd2048;
        rom[2049] = 12'd2049;
        rom[2050] = 12'd2050;
        rom[2051] = 12'd2051;
        rom[2052] = 12'd2052;
        rom[2053] = 12'd2053;
        rom[2054] = 12'd2054;
        rom[2055] = 12'd2055;
        rom[2056] = 12'd2056;
        rom[2057] = 12'd2057;
        rom[2058] = 12'd2058;
        rom[2059] = 12'd2059;
        rom[2060] = 12'd2060;
        rom[2061] = 12'd2061;
        rom[2062] = 12'd2062;
        rom[2063] = 12'd2063;
        rom[2064] = 12'd2064;
        rom[2065] = 12'd2065;
        rom[2066] = 12'd2066;
        rom[2067] = 12'd2067;
        rom[2068] = 12'd2068;
        rom[2069] = 12'd2069;
        rom[2070] = 12'd2070;
        rom[2071] = 12'd2071;
        rom[2072] = 12'd2072;
        rom[2073] = 12'd2073;
        rom[2074] = 12'd2074;
        rom[2075] = 12'd2075;
        rom[2076] = 12'd2076;
        rom[2077] = 12'd2077;
        rom[2078] = 12'd2078;
        rom[2079] = 12'd2079;
        rom[2080] = 12'd2080;
        rom[2081] = 12'd2081;
        rom[2082] = 12'd2082;
        rom[2083] = 12'd2083;
        rom[2084] = 12'd2084;
        rom[2085] = 12'd2085;
        rom[2086] = 12'd2086;
        rom[2087] = 12'd2087;
        rom[2088] = 12'd2088;
        rom[2089] = 12'd2089;
        rom[2090] = 12'd2090;
        rom[2091] = 12'd2091;
        rom[2092] = 12'd2092;
        rom[2093] = 12'd2093;
        rom[2094] = 12'd2094;
        rom[2095] = 12'd2095;
        rom[2096] = 12'd2096;
        rom[2097] = 12'd2097;
        rom[2098] = 12'd2098;
        rom[2099] = 12'd2099;
        rom[2100] = 12'd2100;
        rom[2101] = 12'd2101;
        rom[2102] = 12'd2102;
        rom[2103] = 12'd2103;
        rom[2104] = 12'd2104;
        rom[2105] = 12'd2105;
        rom[2106] = 12'd2106;
        rom[2107] = 12'd2107;
        rom[2108] = 12'd2108;
        rom[2109] = 12'd2109;
        rom[2110] = 12'd2110;
        rom[2111] = 12'd2111;
        rom[2112] = 12'd2112;
        rom[2113] = 12'd2113;
        rom[2114] = 12'd2114;
        rom[2115] = 12'd2115;
        rom[2116] = 12'd2116;
        rom[2117] = 12'd2117;
        rom[2118] = 12'd2118;
        rom[2119] = 12'd2119;
        rom[2120] = 12'd2120;
        rom[2121] = 12'd2121;
        rom[2122] = 12'd2122;
        rom[2123] = 12'd2123;
        rom[2124] = 12'd2124;
        rom[2125] = 12'd2125;
        rom[2126] = 12'd2126;
        rom[2127] = 12'd2127;
        rom[2128] = 12'd2128;
        rom[2129] = 12'd2129;
        rom[2130] = 12'd2130;
        rom[2131] = 12'd2131;
        rom[2132] = 12'd2132;
        rom[2133] = 12'd2133;
        rom[2134] = 12'd2134;
        rom[2135] = 12'd2135;
        rom[2136] = 12'd2136;
        rom[2137] = 12'd2137;
        rom[2138] = 12'd2138;
        rom[2139] = 12'd2139;
        rom[2140] = 12'd2140;
        rom[2141] = 12'd2141;
        rom[2142] = 12'd2142;
        rom[2143] = 12'd2143;
        rom[2144] = 12'd2144;
        rom[2145] = 12'd2145;
        rom[2146] = 12'd2146;
        rom[2147] = 12'd2147;
        rom[2148] = 12'd2148;
        rom[2149] = 12'd2149;
        rom[2150] = 12'd2150;
        rom[2151] = 12'd2151;
        rom[2152] = 12'd2152;
        rom[2153] = 12'd2153;
        rom[2154] = 12'd2154;
        rom[2155] = 12'd2155;
        rom[2156] = 12'd2156;
        rom[2157] = 12'd2157;
        rom[2158] = 12'd2158;
        rom[2159] = 12'd2159;
        rom[2160] = 12'd2160;
        rom[2161] = 12'd2161;
        rom[2162] = 12'd2162;
        rom[2163] = 12'd2163;
        rom[2164] = 12'd2164;
        rom[2165] = 12'd2165;
        rom[2166] = 12'd2166;
        rom[2167] = 12'd2167;
        rom[2168] = 12'd2168;
        rom[2169] = 12'd2169;
        rom[2170] = 12'd2170;
        rom[2171] = 12'd2171;
        rom[2172] = 12'd2172;
        rom[2173] = 12'd2173;
        rom[2174] = 12'd2174;
        rom[2175] = 12'd2175;
        rom[2176] = 12'd2176;
        rom[2177] = 12'd2177;
        rom[2178] = 12'd2178;
        rom[2179] = 12'd2179;
        rom[2180] = 12'd2180;
        rom[2181] = 12'd2181;
        rom[2182] = 12'd2182;
        rom[2183] = 12'd2183;
        rom[2184] = 12'd2184;
        rom[2185] = 12'd2185;
        rom[2186] = 12'd2186;
        rom[2187] = 12'd2187;
        rom[2188] = 12'd2188;
        rom[2189] = 12'd2189;
        rom[2190] = 12'd2190;
        rom[2191] = 12'd2191;
        rom[2192] = 12'd2192;
        rom[2193] = 12'd2193;
        rom[2194] = 12'd2194;
        rom[2195] = 12'd2195;
        rom[2196] = 12'd2196;
        rom[2197] = 12'd2197;
        rom[2198] = 12'd2198;
        rom[2199] = 12'd2199;
        rom[2200] = 12'd2200;
        rom[2201] = 12'd2201;
        rom[2202] = 12'd2202;
        rom[2203] = 12'd2203;
        rom[2204] = 12'd2204;
        rom[2205] = 12'd2205;
        rom[2206] = 12'd2206;
        rom[2207] = 12'd2207;
        rom[2208] = 12'd2208;
        rom[2209] = 12'd2209;
        rom[2210] = 12'd2210;
        rom[2211] = 12'd2211;
        rom[2212] = 12'd2212;
        rom[2213] = 12'd2213;
        rom[2214] = 12'd2214;
        rom[2215] = 12'd2215;
        rom[2216] = 12'd2216;
        rom[2217] = 12'd2217;
        rom[2218] = 12'd2218;
        rom[2219] = 12'd2219;
        rom[2220] = 12'd2220;
        rom[2221] = 12'd2221;
        rom[2222] = 12'd2222;
        rom[2223] = 12'd2223;
        rom[2224] = 12'd2224;
        rom[2225] = 12'd2225;
        rom[2226] = 12'd2226;
        rom[2227] = 12'd2227;
        rom[2228] = 12'd2228;
        rom[2229] = 12'd2229;
        rom[2230] = 12'd2230;
        rom[2231] = 12'd2231;
        rom[2232] = 12'd2232;
        rom[2233] = 12'd2233;
        rom[2234] = 12'd2234;
        rom[2235] = 12'd2235;
        rom[2236] = 12'd2236;
        rom[2237] = 12'd2237;
        rom[2238] = 12'd2238;
        rom[2239] = 12'd2239;
        rom[2240] = 12'd2240;
        rom[2241] = 12'd2241;
        rom[2242] = 12'd2242;
        rom[2243] = 12'd2243;
        rom[2244] = 12'd2244;
        rom[2245] = 12'd2245;
        rom[2246] = 12'd2246;
        rom[2247] = 12'd2247;
        rom[2248] = 12'd2248;
        rom[2249] = 12'd2249;
        rom[2250] = 12'd2250;
        rom[2251] = 12'd2251;
        rom[2252] = 12'd2252;
        rom[2253] = 12'd2253;
        rom[2254] = 12'd2254;
        rom[2255] = 12'd2255;
        rom[2256] = 12'd2256;
        rom[2257] = 12'd2257;
        rom[2258] = 12'd2258;
        rom[2259] = 12'd2259;
        rom[2260] = 12'd2260;
        rom[2261] = 12'd2261;
        rom[2262] = 12'd2262;
        rom[2263] = 12'd2263;
        rom[2264] = 12'd2264;
        rom[2265] = 12'd2265;
        rom[2266] = 12'd2266;
        rom[2267] = 12'd2267;
        rom[2268] = 12'd2268;
        rom[2269] = 12'd2269;
        rom[2270] = 12'd2270;
        rom[2271] = 12'd2271;
        rom[2272] = 12'd2272;
        rom[2273] = 12'd2273;
        rom[2274] = 12'd2274;
        rom[2275] = 12'd2275;
        rom[2276] = 12'd2276;
        rom[2277] = 12'd2277;
        rom[2278] = 12'd2278;
        rom[2279] = 12'd2279;
        rom[2280] = 12'd2280;
        rom[2281] = 12'd2281;
        rom[2282] = 12'd2282;
        rom[2283] = 12'd2283;
        rom[2284] = 12'd2284;
        rom[2285] = 12'd2285;
        rom[2286] = 12'd2286;
        rom[2287] = 12'd2287;
        rom[2288] = 12'd2288;
        rom[2289] = 12'd2289;
        rom[2290] = 12'd2290;
        rom[2291] = 12'd2291;
        rom[2292] = 12'd2292;
        rom[2293] = 12'd2293;
        rom[2294] = 12'd2294;
        rom[2295] = 12'd2295;
        rom[2296] = 12'd2296;
        rom[2297] = 12'd2297;
        rom[2298] = 12'd2298;
        rom[2299] = 12'd2299;
        rom[2300] = 12'd2300;
        rom[2301] = 12'd2301;
        rom[2302] = 12'd2302;
        rom[2303] = 12'd2303;
        rom[2304] = 12'd2304;
        rom[2305] = 12'd2305;
        rom[2306] = 12'd2306;
        rom[2307] = 12'd2307;
        rom[2308] = 12'd2308;
        rom[2309] = 12'd2309;
        rom[2310] = 12'd2310;
        rom[2311] = 12'd2311;
        rom[2312] = 12'd2312;
        rom[2313] = 12'd2313;
        rom[2314] = 12'd2314;
        rom[2315] = 12'd2315;
        rom[2316] = 12'd2316;
        rom[2317] = 12'd2317;
        rom[2318] = 12'd2318;
        rom[2319] = 12'd2319;
        rom[2320] = 12'd2320;
        rom[2321] = 12'd2321;
        rom[2322] = 12'd2322;
        rom[2323] = 12'd2323;
        rom[2324] = 12'd2324;
        rom[2325] = 12'd2325;
        rom[2326] = 12'd2326;
        rom[2327] = 12'd2327;
        rom[2328] = 12'd2328;
        rom[2329] = 12'd2329;
        rom[2330] = 12'd2330;
        rom[2331] = 12'd2331;
        rom[2332] = 12'd2332;
        rom[2333] = 12'd2333;
        rom[2334] = 12'd2334;
        rom[2335] = 12'd2335;
        rom[2336] = 12'd2336;
        rom[2337] = 12'd2337;
        rom[2338] = 12'd2338;
        rom[2339] = 12'd2339;
        rom[2340] = 12'd2340;
        rom[2341] = 12'd2341;
        rom[2342] = 12'd2342;
        rom[2343] = 12'd2343;
        rom[2344] = 12'd2344;
        rom[2345] = 12'd2345;
        rom[2346] = 12'd2346;
        rom[2347] = 12'd2347;
        rom[2348] = 12'd2348;
        rom[2349] = 12'd2349;
        rom[2350] = 12'd2350;
        rom[2351] = 12'd2351;
        rom[2352] = 12'd2352;
        rom[2353] = 12'd2353;
        rom[2354] = 12'd2354;
        rom[2355] = 12'd2355;
        rom[2356] = 12'd2356;
        rom[2357] = 12'd2357;
        rom[2358] = 12'd2358;
        rom[2359] = 12'd2359;
        rom[2360] = 12'd2360;
        rom[2361] = 12'd2361;
        rom[2362] = 12'd2362;
        rom[2363] = 12'd2363;
        rom[2364] = 12'd2364;
        rom[2365] = 12'd2365;
        rom[2366] = 12'd2366;
        rom[2367] = 12'd2367;
        rom[2368] = 12'd2368;
        rom[2369] = 12'd2369;
        rom[2370] = 12'd2370;
        rom[2371] = 12'd2371;
        rom[2372] = 12'd2372;
        rom[2373] = 12'd2373;
        rom[2374] = 12'd2374;
        rom[2375] = 12'd2375;
        rom[2376] = 12'd2376;
        rom[2377] = 12'd2377;
        rom[2378] = 12'd2378;
        rom[2379] = 12'd2379;
        rom[2380] = 12'd2380;
        rom[2381] = 12'd2381;
        rom[2382] = 12'd2382;
        rom[2383] = 12'd2383;
        rom[2384] = 12'd2384;
        rom[2385] = 12'd2385;
        rom[2386] = 12'd2386;
        rom[2387] = 12'd2387;
        rom[2388] = 12'd2388;
        rom[2389] = 12'd2389;
        rom[2390] = 12'd2390;
        rom[2391] = 12'd2391;
        rom[2392] = 12'd2392;
        rom[2393] = 12'd2393;
        rom[2394] = 12'd2394;
        rom[2395] = 12'd2395;
        rom[2396] = 12'd2396;
        rom[2397] = 12'd2397;
        rom[2398] = 12'd2398;
        rom[2399] = 12'd2399;
        rom[2400] = 12'd2400;
        rom[2401] = 12'd2401;
        rom[2402] = 12'd2402;
        rom[2403] = 12'd2403;
        rom[2404] = 12'd2404;
        rom[2405] = 12'd2405;
        rom[2406] = 12'd2406;
        rom[2407] = 12'd2407;
        rom[2408] = 12'd2408;
        rom[2409] = 12'd2409;
        rom[2410] = 12'd2410;
        rom[2411] = 12'd2411;
        rom[2412] = 12'd2412;
        rom[2413] = 12'd2413;
        rom[2414] = 12'd2414;
        rom[2415] = 12'd2415;
        rom[2416] = 12'd2416;
        rom[2417] = 12'd2417;
        rom[2418] = 12'd2418;
        rom[2419] = 12'd2419;
        rom[2420] = 12'd2420;
        rom[2421] = 12'd2421;
        rom[2422] = 12'd2422;
        rom[2423] = 12'd2423;
        rom[2424] = 12'd2424;
        rom[2425] = 12'd2425;
        rom[2426] = 12'd2426;
        rom[2427] = 12'd2427;
        rom[2428] = 12'd2428;
        rom[2429] = 12'd2429;
        rom[2430] = 12'd2430;
        rom[2431] = 12'd2431;
        rom[2432] = 12'd2432;
        rom[2433] = 12'd2433;
        rom[2434] = 12'd2434;
        rom[2435] = 12'd2435;
        rom[2436] = 12'd2436;
        rom[2437] = 12'd2437;
        rom[2438] = 12'd2438;
        rom[2439] = 12'd2439;
        rom[2440] = 12'd2440;
        rom[2441] = 12'd2441;
        rom[2442] = 12'd2442;
        rom[2443] = 12'd2443;
        rom[2444] = 12'd2444;
        rom[2445] = 12'd2445;
        rom[2446] = 12'd2446;
        rom[2447] = 12'd2447;
        rom[2448] = 12'd2448;
        rom[2449] = 12'd2449;
        rom[2450] = 12'd2450;
        rom[2451] = 12'd2451;
        rom[2452] = 12'd2452;
        rom[2453] = 12'd2453;
        rom[2454] = 12'd2454;
        rom[2455] = 12'd2455;
        rom[2456] = 12'd2456;
        rom[2457] = 12'd2457;
        rom[2458] = 12'd2458;
        rom[2459] = 12'd2459;
        rom[2460] = 12'd2460;
        rom[2461] = 12'd2461;
        rom[2462] = 12'd2462;
        rom[2463] = 12'd2463;
        rom[2464] = 12'd2464;
        rom[2465] = 12'd2465;
        rom[2466] = 12'd2466;
        rom[2467] = 12'd2467;
        rom[2468] = 12'd2468;
        rom[2469] = 12'd2469;
        rom[2470] = 12'd2470;
        rom[2471] = 12'd2471;
        rom[2472] = 12'd2472;
        rom[2473] = 12'd2473;
        rom[2474] = 12'd2474;
        rom[2475] = 12'd2475;
        rom[2476] = 12'd2476;
        rom[2477] = 12'd2477;
        rom[2478] = 12'd2478;
        rom[2479] = 12'd2479;
        rom[2480] = 12'd2480;
        rom[2481] = 12'd2481;
        rom[2482] = 12'd2482;
        rom[2483] = 12'd2483;
        rom[2484] = 12'd2484;
        rom[2485] = 12'd2485;
        rom[2486] = 12'd2486;
        rom[2487] = 12'd2487;
        rom[2488] = 12'd2488;
        rom[2489] = 12'd2489;
        rom[2490] = 12'd2490;
        rom[2491] = 12'd2491;
        rom[2492] = 12'd2492;
        rom[2493] = 12'd2493;
        rom[2494] = 12'd2494;
        rom[2495] = 12'd2495;
        rom[2496] = 12'd2496;
        rom[2497] = 12'd2497;
        rom[2498] = 12'd2498;
        rom[2499] = 12'd2499;
        rom[2500] = 12'd2500;
        rom[2501] = 12'd2501;
        rom[2502] = 12'd2502;
        rom[2503] = 12'd2503;
        rom[2504] = 12'd2504;
        rom[2505] = 12'd2505;
        rom[2506] = 12'd2506;
        rom[2507] = 12'd2507;
        rom[2508] = 12'd2508;
        rom[2509] = 12'd2509;
        rom[2510] = 12'd2510;
        rom[2511] = 12'd2511;
        rom[2512] = 12'd2512;
        rom[2513] = 12'd2513;
        rom[2514] = 12'd2514;
        rom[2515] = 12'd2515;
        rom[2516] = 12'd2516;
        rom[2517] = 12'd2517;
        rom[2518] = 12'd2518;
        rom[2519] = 12'd2519;
        rom[2520] = 12'd2520;
        rom[2521] = 12'd2521;
        rom[2522] = 12'd2522;
        rom[2523] = 12'd2523;
        rom[2524] = 12'd2524;
        rom[2525] = 12'd2525;
        rom[2526] = 12'd2526;
        rom[2527] = 12'd2527;
        rom[2528] = 12'd2528;
        rom[2529] = 12'd2529;
        rom[2530] = 12'd2530;
        rom[2531] = 12'd2531;
        rom[2532] = 12'd2532;
        rom[2533] = 12'd2533;
        rom[2534] = 12'd2534;
        rom[2535] = 12'd2535;
        rom[2536] = 12'd2536;
        rom[2537] = 12'd2537;
        rom[2538] = 12'd2538;
        rom[2539] = 12'd2539;
        rom[2540] = 12'd2540;
        rom[2541] = 12'd2541;
        rom[2542] = 12'd2542;
        rom[2543] = 12'd2543;
        rom[2544] = 12'd2544;
        rom[2545] = 12'd2545;
        rom[2546] = 12'd2546;
        rom[2547] = 12'd2547;
        rom[2548] = 12'd2548;
        rom[2549] = 12'd2549;
        rom[2550] = 12'd2550;
        rom[2551] = 12'd2551;
        rom[2552] = 12'd2552;
        rom[2553] = 12'd2553;
        rom[2554] = 12'd2554;
        rom[2555] = 12'd2555;
        rom[2556] = 12'd2556;
        rom[2557] = 12'd2557;
        rom[2558] = 12'd2558;
        rom[2559] = 12'd2559;
        rom[2560] = 12'd2560;
        rom[2561] = 12'd2561;
        rom[2562] = 12'd2562;
        rom[2563] = 12'd2563;
        rom[2564] = 12'd2564;
        rom[2565] = 12'd2565;
        rom[2566] = 12'd2566;
        rom[2567] = 12'd2567;
        rom[2568] = 12'd2568;
        rom[2569] = 12'd2569;
        rom[2570] = 12'd2570;
        rom[2571] = 12'd2571;
        rom[2572] = 12'd2572;
        rom[2573] = 12'd2573;
        rom[2574] = 12'd2574;
        rom[2575] = 12'd2575;
        rom[2576] = 12'd2576;
        rom[2577] = 12'd2577;
        rom[2578] = 12'd2578;
        rom[2579] = 12'd2579;
        rom[2580] = 12'd2580;
        rom[2581] = 12'd2581;
        rom[2582] = 12'd2582;
        rom[2583] = 12'd2583;
        rom[2584] = 12'd2584;
        rom[2585] = 12'd2585;
        rom[2586] = 12'd2586;
        rom[2587] = 12'd2587;
        rom[2588] = 12'd2588;
        rom[2589] = 12'd2589;
        rom[2590] = 12'd2590;
        rom[2591] = 12'd2591;
        rom[2592] = 12'd2592;
        rom[2593] = 12'd2593;
        rom[2594] = 12'd2594;
        rom[2595] = 12'd2595;
        rom[2596] = 12'd2596;
        rom[2597] = 12'd2597;
        rom[2598] = 12'd2598;
        rom[2599] = 12'd2599;
        rom[2600] = 12'd2600;
        rom[2601] = 12'd2601;
        rom[2602] = 12'd2602;
        rom[2603] = 12'd2603;
        rom[2604] = 12'd2604;
        rom[2605] = 12'd2605;
        rom[2606] = 12'd2606;
        rom[2607] = 12'd2607;
        rom[2608] = 12'd2608;
        rom[2609] = 12'd2609;
        rom[2610] = 12'd2610;
        rom[2611] = 12'd2611;
        rom[2612] = 12'd2612;
        rom[2613] = 12'd2613;
        rom[2614] = 12'd2614;
        rom[2615] = 12'd2615;
        rom[2616] = 12'd2616;
        rom[2617] = 12'd2617;
        rom[2618] = 12'd2618;
        rom[2619] = 12'd2619;
        rom[2620] = 12'd2620;
        rom[2621] = 12'd2621;
        rom[2622] = 12'd2622;
        rom[2623] = 12'd2623;
        rom[2624] = 12'd2624;
        rom[2625] = 12'd2625;
        rom[2626] = 12'd2626;
        rom[2627] = 12'd2627;
        rom[2628] = 12'd2628;
        rom[2629] = 12'd2629;
        rom[2630] = 12'd2630;
        rom[2631] = 12'd2631;
        rom[2632] = 12'd2632;
        rom[2633] = 12'd2633;
        rom[2634] = 12'd2634;
        rom[2635] = 12'd2635;
        rom[2636] = 12'd2636;
        rom[2637] = 12'd2637;
        rom[2638] = 12'd2638;
        rom[2639] = 12'd2639;
        rom[2640] = 12'd2640;
        rom[2641] = 12'd2641;
        rom[2642] = 12'd2642;
        rom[2643] = 12'd2643;
        rom[2644] = 12'd2644;
        rom[2645] = 12'd2645;
        rom[2646] = 12'd2646;
        rom[2647] = 12'd2647;
        rom[2648] = 12'd2648;
        rom[2649] = 12'd2649;
        rom[2650] = 12'd2650;
        rom[2651] = 12'd2651;
        rom[2652] = 12'd2652;
        rom[2653] = 12'd2653;
        rom[2654] = 12'd2654;
        rom[2655] = 12'd2655;
        rom[2656] = 12'd2656;
        rom[2657] = 12'd2657;
        rom[2658] = 12'd2658;
        rom[2659] = 12'd2659;
        rom[2660] = 12'd2660;
        rom[2661] = 12'd2661;
        rom[2662] = 12'd2662;
        rom[2663] = 12'd2663;
        rom[2664] = 12'd2664;
        rom[2665] = 12'd2665;
        rom[2666] = 12'd2666;
        rom[2667] = 12'd2667;
        rom[2668] = 12'd2668;
        rom[2669] = 12'd2669;
        rom[2670] = 12'd2670;
        rom[2671] = 12'd2671;
        rom[2672] = 12'd2672;
        rom[2673] = 12'd2673;
        rom[2674] = 12'd2674;
        rom[2675] = 12'd2675;
        rom[2676] = 12'd2676;
        rom[2677] = 12'd2677;
        rom[2678] = 12'd2678;
        rom[2679] = 12'd2679;
        rom[2680] = 12'd2680;
        rom[2681] = 12'd2681;
        rom[2682] = 12'd2682;
        rom[2683] = 12'd2683;
        rom[2684] = 12'd2684;
        rom[2685] = 12'd2685;
        rom[2686] = 12'd2686;
        rom[2687] = 12'd2687;
        rom[2688] = 12'd2688;
        rom[2689] = 12'd2689;
        rom[2690] = 12'd2690;
        rom[2691] = 12'd2691;
        rom[2692] = 12'd2692;
        rom[2693] = 12'd2693;
        rom[2694] = 12'd2694;
        rom[2695] = 12'd2695;
        rom[2696] = 12'd2696;
        rom[2697] = 12'd2697;
        rom[2698] = 12'd2698;
        rom[2699] = 12'd2699;
        rom[2700] = 12'd2700;
        rom[2701] = 12'd2701;
        rom[2702] = 12'd2702;
        rom[2703] = 12'd2703;
        rom[2704] = 12'd2704;
        rom[2705] = 12'd2705;
        rom[2706] = 12'd2706;
        rom[2707] = 12'd2707;
        rom[2708] = 12'd2708;
        rom[2709] = 12'd2709;
        rom[2710] = 12'd2710;
        rom[2711] = 12'd2711;
        rom[2712] = 12'd2712;
        rom[2713] = 12'd2713;
        rom[2714] = 12'd2714;
        rom[2715] = 12'd2715;
        rom[2716] = 12'd2716;
        rom[2717] = 12'd2717;
        rom[2718] = 12'd2718;
        rom[2719] = 12'd2719;
        rom[2720] = 12'd2720;
        rom[2721] = 12'd2721;
        rom[2722] = 12'd2722;
        rom[2723] = 12'd2723;
        rom[2724] = 12'd2724;
        rom[2725] = 12'd2725;
        rom[2726] = 12'd2726;
        rom[2727] = 12'd2727;
        rom[2728] = 12'd2728;
        rom[2729] = 12'd2729;
        rom[2730] = 12'd2730;
        rom[2731] = 12'd2731;
        rom[2732] = 12'd2732;
        rom[2733] = 12'd2733;
        rom[2734] = 12'd2734;
        rom[2735] = 12'd2735;
        rom[2736] = 12'd2736;
        rom[2737] = 12'd2737;
        rom[2738] = 12'd2738;
        rom[2739] = 12'd2739;
        rom[2740] = 12'd2740;
        rom[2741] = 12'd2741;
        rom[2742] = 12'd2742;
        rom[2743] = 12'd2743;
        rom[2744] = 12'd2744;
        rom[2745] = 12'd2745;
        rom[2746] = 12'd2746;
        rom[2747] = 12'd2747;
        rom[2748] = 12'd2748;
        rom[2749] = 12'd2749;
        rom[2750] = 12'd2750;
        rom[2751] = 12'd2751;
        rom[2752] = 12'd2752;
        rom[2753] = 12'd2753;
        rom[2754] = 12'd2754;
        rom[2755] = 12'd2755;
        rom[2756] = 12'd2756;
        rom[2757] = 12'd2757;
        rom[2758] = 12'd2758;
        rom[2759] = 12'd2759;
        rom[2760] = 12'd2760;
        rom[2761] = 12'd2761;
        rom[2762] = 12'd2762;
        rom[2763] = 12'd2763;
        rom[2764] = 12'd2764;
        rom[2765] = 12'd2765;
        rom[2766] = 12'd2766;
        rom[2767] = 12'd2767;
        rom[2768] = 12'd2768;
        rom[2769] = 12'd2769;
        rom[2770] = 12'd2770;
        rom[2771] = 12'd2771;
        rom[2772] = 12'd2772;
        rom[2773] = 12'd2773;
        rom[2774] = 12'd2774;
        rom[2775] = 12'd2775;
        rom[2776] = 12'd2776;
        rom[2777] = 12'd2777;
        rom[2778] = 12'd2778;
        rom[2779] = 12'd2779;
        rom[2780] = 12'd2780;
        rom[2781] = 12'd2781;
        rom[2782] = 12'd2782;
        rom[2783] = 12'd2783;
        rom[2784] = 12'd2784;
        rom[2785] = 12'd2785;
        rom[2786] = 12'd2786;
        rom[2787] = 12'd2787;
        rom[2788] = 12'd2788;
        rom[2789] = 12'd2789;
        rom[2790] = 12'd2790;
        rom[2791] = 12'd2791;
        rom[2792] = 12'd2792;
        rom[2793] = 12'd2793;
        rom[2794] = 12'd2794;
        rom[2795] = 12'd2795;
        rom[2796] = 12'd2796;
        rom[2797] = 12'd2797;
        rom[2798] = 12'd2798;
        rom[2799] = 12'd2799;
        rom[2800] = 12'd2800;
        rom[2801] = 12'd2801;
        rom[2802] = 12'd2802;
        rom[2803] = 12'd2803;
        rom[2804] = 12'd2804;
        rom[2805] = 12'd2805;
        rom[2806] = 12'd2806;
        rom[2807] = 12'd2807;
        rom[2808] = 12'd2808;
        rom[2809] = 12'd2809;
        rom[2810] = 12'd2810;
        rom[2811] = 12'd2811;
        rom[2812] = 12'd2812;
        rom[2813] = 12'd2813;
        rom[2814] = 12'd2814;
        rom[2815] = 12'd2815;
        rom[2816] = 12'd2816;
        rom[2817] = 12'd2817;
        rom[2818] = 12'd2818;
        rom[2819] = 12'd2819;
        rom[2820] = 12'd2820;
        rom[2821] = 12'd2821;
        rom[2822] = 12'd2822;
        rom[2823] = 12'd2823;
        rom[2824] = 12'd2824;
        rom[2825] = 12'd2825;
        rom[2826] = 12'd2826;
        rom[2827] = 12'd2827;
        rom[2828] = 12'd2828;
        rom[2829] = 12'd2829;
        rom[2830] = 12'd2830;
        rom[2831] = 12'd2831;
        rom[2832] = 12'd2832;
        rom[2833] = 12'd2833;
        rom[2834] = 12'd2834;
        rom[2835] = 12'd2835;
        rom[2836] = 12'd2836;
        rom[2837] = 12'd2837;
        rom[2838] = 12'd2838;
        rom[2839] = 12'd2839;
        rom[2840] = 12'd2840;
        rom[2841] = 12'd2841;
        rom[2842] = 12'd2842;
        rom[2843] = 12'd2843;
        rom[2844] = 12'd2844;
        rom[2845] = 12'd2845;
        rom[2846] = 12'd2846;
        rom[2847] = 12'd2847;
        rom[2848] = 12'd2848;
        rom[2849] = 12'd2849;
        rom[2850] = 12'd2850;
        rom[2851] = 12'd2851;
        rom[2852] = 12'd2852;
        rom[2853] = 12'd2853;
        rom[2854] = 12'd2854;
        rom[2855] = 12'd2855;
        rom[2856] = 12'd2856;
        rom[2857] = 12'd2857;
        rom[2858] = 12'd2858;
        rom[2859] = 12'd2859;
        rom[2860] = 12'd2860;
        rom[2861] = 12'd2861;
        rom[2862] = 12'd2862;
        rom[2863] = 12'd2863;
        rom[2864] = 12'd2864;
        rom[2865] = 12'd2865;
        rom[2866] = 12'd2866;
        rom[2867] = 12'd2867;
        rom[2868] = 12'd2868;
        rom[2869] = 12'd2869;
        rom[2870] = 12'd2870;
        rom[2871] = 12'd2871;
        rom[2872] = 12'd2872;
        rom[2873] = 12'd2873;
        rom[2874] = 12'd2874;
        rom[2875] = 12'd2875;
        rom[2876] = 12'd2876;
        rom[2877] = 12'd2877;
        rom[2878] = 12'd2878;
        rom[2879] = 12'd2879;
        rom[2880] = 12'd2880;
        rom[2881] = 12'd2881;
        rom[2882] = 12'd2882;
        rom[2883] = 12'd2883;
        rom[2884] = 12'd2884;
        rom[2885] = 12'd2885;
        rom[2886] = 12'd2886;
        rom[2887] = 12'd2887;
        rom[2888] = 12'd2888;
        rom[2889] = 12'd2889;
        rom[2890] = 12'd2890;
        rom[2891] = 12'd2891;
        rom[2892] = 12'd2892;
        rom[2893] = 12'd2893;
        rom[2894] = 12'd2894;
        rom[2895] = 12'd2895;
        rom[2896] = 12'd2896;
        rom[2897] = 12'd2897;
        rom[2898] = 12'd2898;
        rom[2899] = 12'd2899;
        rom[2900] = 12'd2900;
        rom[2901] = 12'd2901;
        rom[2902] = 12'd2902;
        rom[2903] = 12'd2903;
        rom[2904] = 12'd2904;
        rom[2905] = 12'd2905;
        rom[2906] = 12'd2906;
        rom[2907] = 12'd2907;
        rom[2908] = 12'd2908;
        rom[2909] = 12'd2909;
        rom[2910] = 12'd2910;
        rom[2911] = 12'd2911;
        rom[2912] = 12'd2912;
        rom[2913] = 12'd2913;
        rom[2914] = 12'd2914;
        rom[2915] = 12'd2915;
        rom[2916] = 12'd2916;
        rom[2917] = 12'd2917;
        rom[2918] = 12'd2918;
        rom[2919] = 12'd2919;
        rom[2920] = 12'd2920;
        rom[2921] = 12'd2921;
        rom[2922] = 12'd2922;
        rom[2923] = 12'd2923;
        rom[2924] = 12'd2924;
        rom[2925] = 12'd2925;
        rom[2926] = 12'd2926;
        rom[2927] = 12'd2927;
        rom[2928] = 12'd2928;
        rom[2929] = 12'd2929;
        rom[2930] = 12'd2930;
        rom[2931] = 12'd2931;
        rom[2932] = 12'd2932;
        rom[2933] = 12'd2933;
        rom[2934] = 12'd2934;
        rom[2935] = 12'd2935;
        rom[2936] = 12'd2936;
        rom[2937] = 12'd2937;
        rom[2938] = 12'd2938;
        rom[2939] = 12'd2939;
        rom[2940] = 12'd2940;
        rom[2941] = 12'd2941;
        rom[2942] = 12'd2942;
        rom[2943] = 12'd2943;
        rom[2944] = 12'd2944;
        rom[2945] = 12'd2945;
        rom[2946] = 12'd2946;
        rom[2947] = 12'd2947;
        rom[2948] = 12'd2948;
        rom[2949] = 12'd2949;
        rom[2950] = 12'd2950;
        rom[2951] = 12'd2951;
        rom[2952] = 12'd2952;
        rom[2953] = 12'd2953;
        rom[2954] = 12'd2954;
        rom[2955] = 12'd2955;
        rom[2956] = 12'd2956;
        rom[2957] = 12'd2957;
        rom[2958] = 12'd2958;
        rom[2959] = 12'd2959;
        rom[2960] = 12'd2960;
        rom[2961] = 12'd2961;
        rom[2962] = 12'd2962;
        rom[2963] = 12'd2963;
        rom[2964] = 12'd2964;
        rom[2965] = 12'd2965;
        rom[2966] = 12'd2966;
        rom[2967] = 12'd2967;
        rom[2968] = 12'd2968;
        rom[2969] = 12'd2969;
        rom[2970] = 12'd2970;
        rom[2971] = 12'd2971;
        rom[2972] = 12'd2972;
        rom[2973] = 12'd2973;
        rom[2974] = 12'd2974;
        rom[2975] = 12'd2975;
        rom[2976] = 12'd2976;
        rom[2977] = 12'd2977;
        rom[2978] = 12'd2978;
        rom[2979] = 12'd2979;
        rom[2980] = 12'd2980;
        rom[2981] = 12'd2981;
        rom[2982] = 12'd2982;
        rom[2983] = 12'd2983;
        rom[2984] = 12'd2984;
        rom[2985] = 12'd2985;
        rom[2986] = 12'd2986;
        rom[2987] = 12'd2987;
        rom[2988] = 12'd2988;
        rom[2989] = 12'd2989;
        rom[2990] = 12'd2990;
        rom[2991] = 12'd2991;
        rom[2992] = 12'd2992;
        rom[2993] = 12'd2993;
        rom[2994] = 12'd2994;
        rom[2995] = 12'd2995;
        rom[2996] = 12'd2996;
        rom[2997] = 12'd2997;
        rom[2998] = 12'd2998;
        rom[2999] = 12'd2999;
        rom[3000] = 12'd3000;
        rom[3001] = 12'd3001;
        rom[3002] = 12'd3002;
        rom[3003] = 12'd3003;
        rom[3004] = 12'd3004;
        rom[3005] = 12'd3005;
        rom[3006] = 12'd3006;
        rom[3007] = 12'd3007;
        rom[3008] = 12'd3008;
        rom[3009] = 12'd3009;
        rom[3010] = 12'd3010;
        rom[3011] = 12'd3011;
        rom[3012] = 12'd3012;
        rom[3013] = 12'd3013;
        rom[3014] = 12'd3014;
        rom[3015] = 12'd3015;
        rom[3016] = 12'd3016;
        rom[3017] = 12'd3017;
        rom[3018] = 12'd3018;
        rom[3019] = 12'd3019;
        rom[3020] = 12'd3020;
        rom[3021] = 12'd3021;
        rom[3022] = 12'd3022;
        rom[3023] = 12'd3023;
        rom[3024] = 12'd3024;
        rom[3025] = 12'd3025;
        rom[3026] = 12'd3026;
        rom[3027] = 12'd3027;
        rom[3028] = 12'd3028;
        rom[3029] = 12'd3029;
        rom[3030] = 12'd3030;
        rom[3031] = 12'd3031;
        rom[3032] = 12'd3032;
        rom[3033] = 12'd3033;
        rom[3034] = 12'd3034;
        rom[3035] = 12'd3035;
        rom[3036] = 12'd3036;
        rom[3037] = 12'd3037;
        rom[3038] = 12'd3038;
        rom[3039] = 12'd3039;
        rom[3040] = 12'd3040;
        rom[3041] = 12'd3041;
        rom[3042] = 12'd3042;
        rom[3043] = 12'd3043;
        rom[3044] = 12'd3044;
        rom[3045] = 12'd3045;
        rom[3046] = 12'd3046;
        rom[3047] = 12'd3047;
        rom[3048] = 12'd3048;
        rom[3049] = 12'd3049;
        rom[3050] = 12'd3050;
        rom[3051] = 12'd3051;
        rom[3052] = 12'd3052;
        rom[3053] = 12'd3053;
        rom[3054] = 12'd3054;
        rom[3055] = 12'd3055;
        rom[3056] = 12'd3056;
        rom[3057] = 12'd3057;
        rom[3058] = 12'd3058;
        rom[3059] = 12'd3059;
        rom[3060] = 12'd3060;
        rom[3061] = 12'd3061;
        rom[3062] = 12'd3062;
        rom[3063] = 12'd3063;
        rom[3064] = 12'd3064;
        rom[3065] = 12'd3065;
        rom[3066] = 12'd3066;
        rom[3067] = 12'd3067;
        rom[3068] = 12'd3068;
        rom[3069] = 12'd3069;
        rom[3070] = 12'd3070;
        rom[3071] = 12'd3071;
        rom[3072] = 12'd3072;
        rom[3073] = 12'd3073;
        rom[3074] = 12'd3074;
        rom[3075] = 12'd3075;
        rom[3076] = 12'd3076;
        rom[3077] = 12'd3077;
        rom[3078] = 12'd3078;
        rom[3079] = 12'd3079;
        rom[3080] = 12'd3080;
        rom[3081] = 12'd3081;
        rom[3082] = 12'd3082;
        rom[3083] = 12'd3083;
        rom[3084] = 12'd3084;
        rom[3085] = 12'd3085;
        rom[3086] = 12'd3086;
        rom[3087] = 12'd3087;
        rom[3088] = 12'd3088;
        rom[3089] = 12'd3089;
        rom[3090] = 12'd3090;
        rom[3091] = 12'd3091;
        rom[3092] = 12'd3092;
        rom[3093] = 12'd3093;
        rom[3094] = 12'd3094;
        rom[3095] = 12'd3095;
        rom[3096] = 12'd3096;
        rom[3097] = 12'd3097;
        rom[3098] = 12'd3098;
        rom[3099] = 12'd3099;
        rom[3100] = 12'd3100;
        rom[3101] = 12'd3101;
        rom[3102] = 12'd3102;
        rom[3103] = 12'd3103;
        rom[3104] = 12'd3104;
        rom[3105] = 12'd3105;
        rom[3106] = 12'd3106;
        rom[3107] = 12'd3107;
        rom[3108] = 12'd3108;
        rom[3109] = 12'd3109;
        rom[3110] = 12'd3110;
        rom[3111] = 12'd3111;
        rom[3112] = 12'd3112;
        rom[3113] = 12'd3113;
        rom[3114] = 12'd3114;
        rom[3115] = 12'd3115;
        rom[3116] = 12'd3116;
        rom[3117] = 12'd3117;
        rom[3118] = 12'd3118;
        rom[3119] = 12'd3119;
        rom[3120] = 12'd3120;
        rom[3121] = 12'd3121;
        rom[3122] = 12'd3122;
        rom[3123] = 12'd3123;
        rom[3124] = 12'd3124;
        rom[3125] = 12'd3125;
        rom[3126] = 12'd3126;
        rom[3127] = 12'd3127;
        rom[3128] = 12'd3128;
        rom[3129] = 12'd3129;
        rom[3130] = 12'd3130;
        rom[3131] = 12'd3131;
        rom[3132] = 12'd3132;
        rom[3133] = 12'd3133;
        rom[3134] = 12'd3134;
        rom[3135] = 12'd3135;
        rom[3136] = 12'd3136;
        rom[3137] = 12'd3137;
        rom[3138] = 12'd3138;
        rom[3139] = 12'd3139;
        rom[3140] = 12'd3140;
        rom[3141] = 12'd3141;
        rom[3142] = 12'd3142;
        rom[3143] = 12'd3143;
        rom[3144] = 12'd3144;
        rom[3145] = 12'd3145;
        rom[3146] = 12'd3146;
        rom[3147] = 12'd3147;
        rom[3148] = 12'd3148;
        rom[3149] = 12'd3149;
        rom[3150] = 12'd3150;
        rom[3151] = 12'd3151;
        rom[3152] = 12'd3152;
        rom[3153] = 12'd3153;
        rom[3154] = 12'd3154;
        rom[3155] = 12'd3155;
        rom[3156] = 12'd3156;
        rom[3157] = 12'd3157;
        rom[3158] = 12'd3158;
        rom[3159] = 12'd3159;
        rom[3160] = 12'd3160;
        rom[3161] = 12'd3161;
        rom[3162] = 12'd3162;
        rom[3163] = 12'd3163;
        rom[3164] = 12'd3164;
        rom[3165] = 12'd3165;
        rom[3166] = 12'd3166;
        rom[3167] = 12'd3167;
        rom[3168] = 12'd3168;
        rom[3169] = 12'd3169;
        rom[3170] = 12'd3170;
        rom[3171] = 12'd3171;
        rom[3172] = 12'd3172;
        rom[3173] = 12'd3173;
        rom[3174] = 12'd3174;
        rom[3175] = 12'd3175;
        rom[3176] = 12'd3176;
        rom[3177] = 12'd3177;
        rom[3178] = 12'd3178;
        rom[3179] = 12'd3179;
        rom[3180] = 12'd3180;
        rom[3181] = 12'd3181;
        rom[3182] = 12'd3182;
        rom[3183] = 12'd3183;
        rom[3184] = 12'd3184;
        rom[3185] = 12'd3185;
        rom[3186] = 12'd3186;
        rom[3187] = 12'd3187;
        rom[3188] = 12'd3188;
        rom[3189] = 12'd3189;
        rom[3190] = 12'd3190;
        rom[3191] = 12'd3191;
        rom[3192] = 12'd3192;
        rom[3193] = 12'd3193;
        rom[3194] = 12'd3194;
        rom[3195] = 12'd3195;
        rom[3196] = 12'd3196;
        rom[3197] = 12'd3197;
        rom[3198] = 12'd3198;
        rom[3199] = 12'd3199;
        rom[3200] = 12'd3200;
        rom[3201] = 12'd3201;
        rom[3202] = 12'd3202;
        rom[3203] = 12'd3203;
        rom[3204] = 12'd3204;
        rom[3205] = 12'd3205;
        rom[3206] = 12'd3206;
        rom[3207] = 12'd3207;
        rom[3208] = 12'd3208;
        rom[3209] = 12'd3209;
        rom[3210] = 12'd3210;
        rom[3211] = 12'd3211;
        rom[3212] = 12'd3212;
        rom[3213] = 12'd3213;
        rom[3214] = 12'd3214;
        rom[3215] = 12'd3215;
        rom[3216] = 12'd3216;
        rom[3217] = 12'd3217;
        rom[3218] = 12'd3218;
        rom[3219] = 12'd3219;
        rom[3220] = 12'd3220;
        rom[3221] = 12'd3221;
        rom[3222] = 12'd3222;
        rom[3223] = 12'd3223;
        rom[3224] = 12'd3224;
        rom[3225] = 12'd3225;
        rom[3226] = 12'd3226;
        rom[3227] = 12'd3227;
        rom[3228] = 12'd3228;
        rom[3229] = 12'd3229;
        rom[3230] = 12'd3230;
        rom[3231] = 12'd3231;
        rom[3232] = 12'd3232;
        rom[3233] = 12'd3233;
        rom[3234] = 12'd3234;
        rom[3235] = 12'd3235;
        rom[3236] = 12'd3236;
        rom[3237] = 12'd3237;
        rom[3238] = 12'd3238;
        rom[3239] = 12'd3239;
        rom[3240] = 12'd3240;
        rom[3241] = 12'd3241;
        rom[3242] = 12'd3242;
        rom[3243] = 12'd3243;
        rom[3244] = 12'd3244;
        rom[3245] = 12'd3245;
        rom[3246] = 12'd3246;
        rom[3247] = 12'd3247;
        rom[3248] = 12'd3248;
        rom[3249] = 12'd3249;
        rom[3250] = 12'd3250;
        rom[3251] = 12'd3251;
        rom[3252] = 12'd3252;
        rom[3253] = 12'd3253;
        rom[3254] = 12'd3254;
        rom[3255] = 12'd3255;
        rom[3256] = 12'd3256;
        rom[3257] = 12'd3257;
        rom[3258] = 12'd3258;
        rom[3259] = 12'd3259;
        rom[3260] = 12'd3260;
        rom[3261] = 12'd3261;
        rom[3262] = 12'd3262;
        rom[3263] = 12'd3263;
        rom[3264] = 12'd3264;
        rom[3265] = 12'd3265;
        rom[3266] = 12'd3266;
        rom[3267] = 12'd3267;
        rom[3268] = 12'd3268;
        rom[3269] = 12'd3269;
        rom[3270] = 12'd3270;
        rom[3271] = 12'd3271;
        rom[3272] = 12'd3272;
        rom[3273] = 12'd3273;
        rom[3274] = 12'd3274;
        rom[3275] = 12'd3275;
        rom[3276] = 12'd3276;
        rom[3277] = 12'd3277;
        rom[3278] = 12'd3278;
        rom[3279] = 12'd3279;
        rom[3280] = 12'd3280;
        rom[3281] = 12'd3281;
        rom[3282] = 12'd3282;
        rom[3283] = 12'd3283;
        rom[3284] = 12'd3284;
        rom[3285] = 12'd3285;
        rom[3286] = 12'd3286;
        rom[3287] = 12'd3287;
        rom[3288] = 12'd3288;
        rom[3289] = 12'd3289;
        rom[3290] = 12'd3290;
        rom[3291] = 12'd3291;
        rom[3292] = 12'd3292;
        rom[3293] = 12'd3293;
        rom[3294] = 12'd3294;
        rom[3295] = 12'd3295;
        rom[3296] = 12'd3296;
        rom[3297] = 12'd3297;
        rom[3298] = 12'd3298;
        rom[3299] = 12'd3299;
        rom[3300] = 12'd3300;
        rom[3301] = 12'd3301;
        rom[3302] = 12'd3302;
        rom[3303] = 12'd3303;
        rom[3304] = 12'd3304;
        rom[3305] = 12'd3305;
        rom[3306] = 12'd3306;
        rom[3307] = 12'd3307;
        rom[3308] = 12'd3308;
        rom[3309] = 12'd3309;
        rom[3310] = 12'd3310;
        rom[3311] = 12'd3311;
        rom[3312] = 12'd3312;
        rom[3313] = 12'd3313;
        rom[3314] = 12'd3314;
        rom[3315] = 12'd3315;
        rom[3316] = 12'd3316;
        rom[3317] = 12'd3317;
        rom[3318] = 12'd3318;
        rom[3319] = 12'd3319;
        rom[3320] = 12'd3320;
        rom[3321] = 12'd3321;
        rom[3322] = 12'd3322;
        rom[3323] = 12'd3323;
        rom[3324] = 12'd3324;
        rom[3325] = 12'd3325;
        rom[3326] = 12'd3326;
        rom[3327] = 12'd3327;
        rom[3328] = 12'd3328;
        rom[3329] = 12'd3329;
        rom[3330] = 12'd3330;
        rom[3331] = 12'd3331;
        rom[3332] = 12'd3332;
        rom[3333] = 12'd3333;
        rom[3334] = 12'd3334;
        rom[3335] = 12'd3335;
        rom[3336] = 12'd3336;
        rom[3337] = 12'd3337;
        rom[3338] = 12'd3338;
        rom[3339] = 12'd3339;
        rom[3340] = 12'd3340;
        rom[3341] = 12'd3341;
        rom[3342] = 12'd3342;
        rom[3343] = 12'd3343;
        rom[3344] = 12'd3344;
        rom[3345] = 12'd3345;
        rom[3346] = 12'd3346;
        rom[3347] = 12'd3347;
        rom[3348] = 12'd3348;
        rom[3349] = 12'd3349;
        rom[3350] = 12'd3350;
        rom[3351] = 12'd3351;
        rom[3352] = 12'd3352;
        rom[3353] = 12'd3353;
        rom[3354] = 12'd3354;
        rom[3355] = 12'd3355;
        rom[3356] = 12'd3356;
        rom[3357] = 12'd3357;
        rom[3358] = 12'd3358;
        rom[3359] = 12'd3359;
        rom[3360] = 12'd3360;
        rom[3361] = 12'd3361;
        rom[3362] = 12'd3362;
        rom[3363] = 12'd3363;
        rom[3364] = 12'd3364;
        rom[3365] = 12'd3365;
        rom[3366] = 12'd3366;
        rom[3367] = 12'd3367;
        rom[3368] = 12'd3368;
        rom[3369] = 12'd3369;
        rom[3370] = 12'd3370;
        rom[3371] = 12'd3371;
        rom[3372] = 12'd3372;
        rom[3373] = 12'd3373;
        rom[3374] = 12'd3374;
        rom[3375] = 12'd3375;
        rom[3376] = 12'd3376;
        rom[3377] = 12'd3377;
        rom[3378] = 12'd3378;
        rom[3379] = 12'd3379;
        rom[3380] = 12'd3380;
        rom[3381] = 12'd3381;
        rom[3382] = 12'd3382;
        rom[3383] = 12'd3383;
        rom[3384] = 12'd3384;
        rom[3385] = 12'd3385;
        rom[3386] = 12'd3386;
        rom[3387] = 12'd3387;
        rom[3388] = 12'd3388;
        rom[3389] = 12'd3389;
        rom[3390] = 12'd3390;
        rom[3391] = 12'd3391;
        rom[3392] = 12'd3392;
        rom[3393] = 12'd3393;
        rom[3394] = 12'd3394;
        rom[3395] = 12'd3395;
        rom[3396] = 12'd3396;
        rom[3397] = 12'd3397;
        rom[3398] = 12'd3398;
        rom[3399] = 12'd3399;
        rom[3400] = 12'd3400;
        rom[3401] = 12'd3401;
        rom[3402] = 12'd3402;
        rom[3403] = 12'd3403;
        rom[3404] = 12'd3404;
        rom[3405] = 12'd3405;
        rom[3406] = 12'd3406;
        rom[3407] = 12'd3407;
        rom[3408] = 12'd3408;
        rom[3409] = 12'd3409;
        rom[3410] = 12'd3410;
        rom[3411] = 12'd3411;
        rom[3412] = 12'd3412;
        rom[3413] = 12'd3413;
        rom[3414] = 12'd3414;
        rom[3415] = 12'd3415;
        rom[3416] = 12'd3416;
        rom[3417] = 12'd3417;
        rom[3418] = 12'd3418;
        rom[3419] = 12'd3419;
        rom[3420] = 12'd3420;
        rom[3421] = 12'd3421;
        rom[3422] = 12'd3422;
        rom[3423] = 12'd3423;
        rom[3424] = 12'd3424;
        rom[3425] = 12'd3425;
        rom[3426] = 12'd3426;
        rom[3427] = 12'd3427;
        rom[3428] = 12'd3428;
        rom[3429] = 12'd3429;
        rom[3430] = 12'd3430;
        rom[3431] = 12'd3431;
        rom[3432] = 12'd3432;
        rom[3433] = 12'd3433;
        rom[3434] = 12'd3434;
        rom[3435] = 12'd3435;
        rom[3436] = 12'd3436;
        rom[3437] = 12'd3437;
        rom[3438] = 12'd3438;
        rom[3439] = 12'd3439;
        rom[3440] = 12'd3440;
        rom[3441] = 12'd3441;
        rom[3442] = 12'd3442;
        rom[3443] = 12'd3443;
        rom[3444] = 12'd3444;
        rom[3445] = 12'd3445;
        rom[3446] = 12'd3446;
        rom[3447] = 12'd3447;
        rom[3448] = 12'd3448;
        rom[3449] = 12'd3449;
        rom[3450] = 12'd3450;
        rom[3451] = 12'd3451;
        rom[3452] = 12'd3452;
        rom[3453] = 12'd3453;
        rom[3454] = 12'd3454;
        rom[3455] = 12'd3455;
        rom[3456] = 12'd3456;
        rom[3457] = 12'd3457;
        rom[3458] = 12'd3458;
        rom[3459] = 12'd3459;
        rom[3460] = 12'd3460;
        rom[3461] = 12'd3461;
        rom[3462] = 12'd3462;
        rom[3463] = 12'd3463;
        rom[3464] = 12'd3464;
        rom[3465] = 12'd3465;
        rom[3466] = 12'd3466;
        rom[3467] = 12'd3467;
        rom[3468] = 12'd3468;
        rom[3469] = 12'd3469;
        rom[3470] = 12'd3470;
        rom[3471] = 12'd3471;
        rom[3472] = 12'd3472;
        rom[3473] = 12'd3473;
        rom[3474] = 12'd3474;
        rom[3475] = 12'd3475;
        rom[3476] = 12'd3476;
        rom[3477] = 12'd3477;
        rom[3478] = 12'd3478;
        rom[3479] = 12'd3479;
        rom[3480] = 12'd3480;
        rom[3481] = 12'd3481;
        rom[3482] = 12'd3482;
        rom[3483] = 12'd3483;
        rom[3484] = 12'd3484;
        rom[3485] = 12'd3485;
        rom[3486] = 12'd3486;
        rom[3487] = 12'd3487;
        rom[3488] = 12'd3488;
        rom[3489] = 12'd3489;
        rom[3490] = 12'd3490;
        rom[3491] = 12'd3491;
        rom[3492] = 12'd3492;
        rom[3493] = 12'd3493;
        rom[3494] = 12'd3494;
        rom[3495] = 12'd3495;
        rom[3496] = 12'd3496;
        rom[3497] = 12'd3497;
        rom[3498] = 12'd3498;
        rom[3499] = 12'd3499;
        rom[3500] = 12'd3500;
        rom[3501] = 12'd3501;
        rom[3502] = 12'd3502;
        rom[3503] = 12'd3503;
        rom[3504] = 12'd3504;
        rom[3505] = 12'd3505;
        rom[3506] = 12'd3506;
        rom[3507] = 12'd3507;
        rom[3508] = 12'd3508;
        rom[3509] = 12'd3509;
        rom[3510] = 12'd3510;
        rom[3511] = 12'd3511;
        rom[3512] = 12'd3512;
        rom[3513] = 12'd3513;
        rom[3514] = 12'd3514;
        rom[3515] = 12'd3515;
        rom[3516] = 12'd3516;
        rom[3517] = 12'd3517;
        rom[3518] = 12'd3518;
        rom[3519] = 12'd3519;
        rom[3520] = 12'd3520;
        rom[3521] = 12'd3521;
        rom[3522] = 12'd3522;
        rom[3523] = 12'd3523;
        rom[3524] = 12'd3524;
        rom[3525] = 12'd3525;
        rom[3526] = 12'd3526;
        rom[3527] = 12'd3527;
        rom[3528] = 12'd3528;
        rom[3529] = 12'd3529;
        rom[3530] = 12'd3530;
        rom[3531] = 12'd3531;
        rom[3532] = 12'd3532;
        rom[3533] = 12'd3533;
        rom[3534] = 12'd3534;
        rom[3535] = 12'd3535;
        rom[3536] = 12'd3536;
        rom[3537] = 12'd3537;
        rom[3538] = 12'd3538;
        rom[3539] = 12'd3539;
        rom[3540] = 12'd3540;
        rom[3541] = 12'd3541;
        rom[3542] = 12'd3542;
        rom[3543] = 12'd3543;
        rom[3544] = 12'd3544;
        rom[3545] = 12'd3545;
        rom[3546] = 12'd3546;
        rom[3547] = 12'd3547;
        rom[3548] = 12'd3548;
        rom[3549] = 12'd3549;
        rom[3550] = 12'd3550;
        rom[3551] = 12'd3551;
        rom[3552] = 12'd3552;
        rom[3553] = 12'd3553;
        rom[3554] = 12'd3554;
        rom[3555] = 12'd3555;
        rom[3556] = 12'd3556;
        rom[3557] = 12'd3557;
        rom[3558] = 12'd3558;
        rom[3559] = 12'd3559;
        rom[3560] = 12'd3560;
        rom[3561] = 12'd3561;
        rom[3562] = 12'd3562;
        rom[3563] = 12'd3563;
        rom[3564] = 12'd3564;
        rom[3565] = 12'd3565;
        rom[3566] = 12'd3566;
        rom[3567] = 12'd3567;
        rom[3568] = 12'd3568;
        rom[3569] = 12'd3569;
        rom[3570] = 12'd3570;
        rom[3571] = 12'd3571;
        rom[3572] = 12'd3572;
        rom[3573] = 12'd3573;
        rom[3574] = 12'd3574;
        rom[3575] = 12'd3575;
        rom[3576] = 12'd3576;
        rom[3577] = 12'd3577;
        rom[3578] = 12'd3578;
        rom[3579] = 12'd3579;
        rom[3580] = 12'd3580;
        rom[3581] = 12'd3581;
        rom[3582] = 12'd3582;
        rom[3583] = 12'd3583;
        rom[3584] = 12'd3584;
        rom[3585] = 12'd3585;
        rom[3586] = 12'd3586;
        rom[3587] = 12'd3587;
        rom[3588] = 12'd3588;
        rom[3589] = 12'd3589;
        rom[3590] = 12'd3590;
        rom[3591] = 12'd3591;
        rom[3592] = 12'd3592;
        rom[3593] = 12'd3593;
        rom[3594] = 12'd3594;
        rom[3595] = 12'd3595;
        rom[3596] = 12'd3596;
        rom[3597] = 12'd3597;
        rom[3598] = 12'd3598;
        rom[3599] = 12'd3599;
        rom[3600] = 12'd3600;
        rom[3601] = 12'd3601;
        rom[3602] = 12'd3602;
        rom[3603] = 12'd3603;
        rom[3604] = 12'd3604;
        rom[3605] = 12'd3605;
        rom[3606] = 12'd3606;
        rom[3607] = 12'd3607;
        rom[3608] = 12'd3608;
        rom[3609] = 12'd3609;
        rom[3610] = 12'd3610;
        rom[3611] = 12'd3611;
        rom[3612] = 12'd3612;
        rom[3613] = 12'd3613;
        rom[3614] = 12'd3614;
        rom[3615] = 12'd3615;
        rom[3616] = 12'd3616;
        rom[3617] = 12'd3617;
        rom[3618] = 12'd3618;
        rom[3619] = 12'd3619;
        rom[3620] = 12'd3620;
        rom[3621] = 12'd3621;
        rom[3622] = 12'd3622;
        rom[3623] = 12'd3623;
        rom[3624] = 12'd3624;
        rom[3625] = 12'd3625;
        rom[3626] = 12'd3626;
        rom[3627] = 12'd3627;
        rom[3628] = 12'd3628;
        rom[3629] = 12'd3629;
        rom[3630] = 12'd3630;
        rom[3631] = 12'd3631;
        rom[3632] = 12'd3632;
        rom[3633] = 12'd3633;
        rom[3634] = 12'd3634;
        rom[3635] = 12'd3635;
        rom[3636] = 12'd3636;
        rom[3637] = 12'd3637;
        rom[3638] = 12'd3638;
        rom[3639] = 12'd3639;
        rom[3640] = 12'd3640;
        rom[3641] = 12'd3641;
        rom[3642] = 12'd3642;
        rom[3643] = 12'd3643;
        rom[3644] = 12'd3644;
        rom[3645] = 12'd3645;
        rom[3646] = 12'd3646;
        rom[3647] = 12'd3647;
        rom[3648] = 12'd3648;
        rom[3649] = 12'd3649;
        rom[3650] = 12'd3650;
        rom[3651] = 12'd3651;
        rom[3652] = 12'd3652;
        rom[3653] = 12'd3653;
        rom[3654] = 12'd3654;
        rom[3655] = 12'd3655;
        rom[3656] = 12'd3656;
        rom[3657] = 12'd3657;
        rom[3658] = 12'd3658;
        rom[3659] = 12'd3659;
        rom[3660] = 12'd3660;
        rom[3661] = 12'd3661;
        rom[3662] = 12'd3662;
        rom[3663] = 12'd3663;
        rom[3664] = 12'd3664;
        rom[3665] = 12'd3665;
        rom[3666] = 12'd3666;
        rom[3667] = 12'd3667;
        rom[3668] = 12'd3668;
        rom[3669] = 12'd3669;
        rom[3670] = 12'd3670;
        rom[3671] = 12'd3671;
        rom[3672] = 12'd3672;
        rom[3673] = 12'd3673;
        rom[3674] = 12'd3674;
        rom[3675] = 12'd3675;
        rom[3676] = 12'd3676;
        rom[3677] = 12'd3677;
        rom[3678] = 12'd3678;
        rom[3679] = 12'd3679;
        rom[3680] = 12'd3680;
        rom[3681] = 12'd3681;
        rom[3682] = 12'd3682;
        rom[3683] = 12'd3683;
        rom[3684] = 12'd3684;
        rom[3685] = 12'd3685;
        rom[3686] = 12'd3686;
        rom[3687] = 12'd3687;
        rom[3688] = 12'd3688;
        rom[3689] = 12'd3689;
        rom[3690] = 12'd3690;
        rom[3691] = 12'd3691;
        rom[3692] = 12'd3692;
        rom[3693] = 12'd3693;
        rom[3694] = 12'd3694;
        rom[3695] = 12'd3695;
        rom[3696] = 12'd3696;
        rom[3697] = 12'd3697;
        rom[3698] = 12'd3698;
        rom[3699] = 12'd3699;
        rom[3700] = 12'd3700;
        rom[3701] = 12'd3701;
        rom[3702] = 12'd3702;
        rom[3703] = 12'd3703;
        rom[3704] = 12'd3704;
        rom[3705] = 12'd3705;
        rom[3706] = 12'd3706;
        rom[3707] = 12'd3707;
        rom[3708] = 12'd3708;
        rom[3709] = 12'd3709;
        rom[3710] = 12'd3710;
        rom[3711] = 12'd3711;
        rom[3712] = 12'd3712;
        rom[3713] = 12'd3713;
        rom[3714] = 12'd3714;
        rom[3715] = 12'd3715;
        rom[3716] = 12'd3716;
        rom[3717] = 12'd3717;
        rom[3718] = 12'd3718;
        rom[3719] = 12'd3719;
        rom[3720] = 12'd3720;
        rom[3721] = 12'd3721;
        rom[3722] = 12'd3722;
        rom[3723] = 12'd3723;
        rom[3724] = 12'd3724;
        rom[3725] = 12'd3725;
        rom[3726] = 12'd3726;
        rom[3727] = 12'd3727;
        rom[3728] = 12'd3728;
        rom[3729] = 12'd3729;
        rom[3730] = 12'd3730;
        rom[3731] = 12'd3731;
        rom[3732] = 12'd3732;
        rom[3733] = 12'd3733;
        rom[3734] = 12'd3734;
        rom[3735] = 12'd3735;
        rom[3736] = 12'd3736;
        rom[3737] = 12'd3737;
        rom[3738] = 12'd3738;
        rom[3739] = 12'd3739;
        rom[3740] = 12'd3740;
        rom[3741] = 12'd3741;
        rom[3742] = 12'd3742;
        rom[3743] = 12'd3743;
        rom[3744] = 12'd3744;
        rom[3745] = 12'd3745;
        rom[3746] = 12'd3746;
        rom[3747] = 12'd3747;
        rom[3748] = 12'd3748;
        rom[3749] = 12'd3749;
        rom[3750] = 12'd3750;
        rom[3751] = 12'd3751;
        rom[3752] = 12'd3752;
        rom[3753] = 12'd3753;
        rom[3754] = 12'd3754;
        rom[3755] = 12'd3755;
        rom[3756] = 12'd3756;
        rom[3757] = 12'd3757;
        rom[3758] = 12'd3758;
        rom[3759] = 12'd3759;
        rom[3760] = 12'd3760;
        rom[3761] = 12'd3761;
        rom[3762] = 12'd3762;
        rom[3763] = 12'd3763;
        rom[3764] = 12'd3764;
        rom[3765] = 12'd3765;
        rom[3766] = 12'd3766;
        rom[3767] = 12'd3767;
        rom[3768] = 12'd3768;
        rom[3769] = 12'd3769;
        rom[3770] = 12'd3770;
        rom[3771] = 12'd3771;
        rom[3772] = 12'd3772;
        rom[3773] = 12'd3773;
        rom[3774] = 12'd3774;
        rom[3775] = 12'd3775;
        rom[3776] = 12'd3776;
        rom[3777] = 12'd3777;
        rom[3778] = 12'd3778;
        rom[3779] = 12'd3779;
        rom[3780] = 12'd3780;
        rom[3781] = 12'd3781;
        rom[3782] = 12'd3782;
        rom[3783] = 12'd3783;
        rom[3784] = 12'd3784;
        rom[3785] = 12'd3785;
        rom[3786] = 12'd3786;
        rom[3787] = 12'd3787;
        rom[3788] = 12'd3788;
        rom[3789] = 12'd3789;
        rom[3790] = 12'd3790;
        rom[3791] = 12'd3791;
        rom[3792] = 12'd3792;
        rom[3793] = 12'd3793;
        rom[3794] = 12'd3794;
        rom[3795] = 12'd3795;
        rom[3796] = 12'd3796;
        rom[3797] = 12'd3797;
        rom[3798] = 12'd3798;
        rom[3799] = 12'd3799;
        rom[3800] = 12'd3800;
        rom[3801] = 12'd3801;
        rom[3802] = 12'd3802;
        rom[3803] = 12'd3803;
        rom[3804] = 12'd3804;
        rom[3805] = 12'd3805;
        rom[3806] = 12'd3806;
        rom[3807] = 12'd3807;
        rom[3808] = 12'd3808;
        rom[3809] = 12'd3809;
        rom[3810] = 12'd3810;
        rom[3811] = 12'd3811;
        rom[3812] = 12'd3812;
        rom[3813] = 12'd3813;
        rom[3814] = 12'd3814;
        rom[3815] = 12'd3815;
        rom[3816] = 12'd3816;
        rom[3817] = 12'd3817;
        rom[3818] = 12'd3818;
        rom[3819] = 12'd3819;
        rom[3820] = 12'd3820;
        rom[3821] = 12'd3821;
        rom[3822] = 12'd3822;
        rom[3823] = 12'd3823;
        rom[3824] = 12'd3824;
        rom[3825] = 12'd3825;
        rom[3826] = 12'd3826;
        rom[3827] = 12'd3827;
        rom[3828] = 12'd3828;
        rom[3829] = 12'd3829;
        rom[3830] = 12'd3830;
        rom[3831] = 12'd3831;
        rom[3832] = 12'd3832;
        rom[3833] = 12'd3833;
        rom[3834] = 12'd3834;
        rom[3835] = 12'd3835;
        rom[3836] = 12'd3836;
        rom[3837] = 12'd3837;
        rom[3838] = 12'd3838;
        rom[3839] = 12'd3839;
        rom[3840] = 12'd3840;
        rom[3841] = 12'd3841;
        rom[3842] = 12'd3842;
        rom[3843] = 12'd3843;
        rom[3844] = 12'd3844;
        rom[3845] = 12'd3845;
        rom[3846] = 12'd3846;
        rom[3847] = 12'd3847;
        rom[3848] = 12'd3848;
        rom[3849] = 12'd3849;
        rom[3850] = 12'd3850;
        rom[3851] = 12'd3851;
        rom[3852] = 12'd3852;
        rom[3853] = 12'd3853;
        rom[3854] = 12'd3854;
        rom[3855] = 12'd3855;
        rom[3856] = 12'd3856;
        rom[3857] = 12'd3857;
        rom[3858] = 12'd3858;
        rom[3859] = 12'd3859;
        rom[3860] = 12'd3860;
        rom[3861] = 12'd3861;
        rom[3862] = 12'd3862;
        rom[3863] = 12'd3863;
        rom[3864] = 12'd3864;
        rom[3865] = 12'd3865;
        rom[3866] = 12'd3866;
        rom[3867] = 12'd3867;
        rom[3868] = 12'd3868;
        rom[3869] = 12'd3869;
        rom[3870] = 12'd3870;
        rom[3871] = 12'd3871;
        rom[3872] = 12'd3872;
        rom[3873] = 12'd3873;
        rom[3874] = 12'd3874;
        rom[3875] = 12'd3875;
        rom[3876] = 12'd3876;
        rom[3877] = 12'd3877;
        rom[3878] = 12'd3878;
        rom[3879] = 12'd3879;
        rom[3880] = 12'd3880;
        rom[3881] = 12'd3881;
        rom[3882] = 12'd3882;
        rom[3883] = 12'd3883;
        rom[3884] = 12'd3884;
        rom[3885] = 12'd3885;
        rom[3886] = 12'd3886;
        rom[3887] = 12'd3887;
        rom[3888] = 12'd3888;
        rom[3889] = 12'd3889;
        rom[3890] = 12'd3890;
        rom[3891] = 12'd3891;
        rom[3892] = 12'd3892;
        rom[3893] = 12'd3893;
        rom[3894] = 12'd3894;
        rom[3895] = 12'd3895;
        rom[3896] = 12'd3896;
        rom[3897] = 12'd3897;
        rom[3898] = 12'd3898;
        rom[3899] = 12'd3899;
        rom[3900] = 12'd3900;
        rom[3901] = 12'd3901;
        rom[3902] = 12'd3902;
        rom[3903] = 12'd3903;
        rom[3904] = 12'd3904;
        rom[3905] = 12'd3905;
        rom[3906] = 12'd3906;
        rom[3907] = 12'd3907;
        rom[3908] = 12'd3908;
        rom[3909] = 12'd3909;
        rom[3910] = 12'd3910;
        rom[3911] = 12'd3911;
        rom[3912] = 12'd3912;
        rom[3913] = 12'd3913;
        rom[3914] = 12'd3914;
        rom[3915] = 12'd3915;
        rom[3916] = 12'd3916;
        rom[3917] = 12'd3917;
        rom[3918] = 12'd3918;
        rom[3919] = 12'd3919;
        rom[3920] = 12'd3920;
        rom[3921] = 12'd3921;
        rom[3922] = 12'd3922;
        rom[3923] = 12'd3923;
        rom[3924] = 12'd3924;
        rom[3925] = 12'd3925;
        rom[3926] = 12'd3926;
        rom[3927] = 12'd3927;
        rom[3928] = 12'd3928;
        rom[3929] = 12'd3929;
        rom[3930] = 12'd3930;
        rom[3931] = 12'd3931;
        rom[3932] = 12'd3932;
        rom[3933] = 12'd3933;
        rom[3934] = 12'd3934;
        rom[3935] = 12'd3935;
        rom[3936] = 12'd3936;
        rom[3937] = 12'd3937;
        rom[3938] = 12'd3938;
        rom[3939] = 12'd3939;
        rom[3940] = 12'd3940;
        rom[3941] = 12'd3941;
        rom[3942] = 12'd3942;
        rom[3943] = 12'd3943;
        rom[3944] = 12'd3944;
        rom[3945] = 12'd3945;
        rom[3946] = 12'd3946;
        rom[3947] = 12'd3947;
        rom[3948] = 12'd3948;
        rom[3949] = 12'd3949;
        rom[3950] = 12'd3950;
        rom[3951] = 12'd3951;
        rom[3952] = 12'd3952;
        rom[3953] = 12'd3953;
        rom[3954] = 12'd3954;
        rom[3955] = 12'd3955;
        rom[3956] = 12'd3956;
        rom[3957] = 12'd3957;
        rom[3958] = 12'd3958;
        rom[3959] = 12'd3959;
        rom[3960] = 12'd3960;
        rom[3961] = 12'd3961;
        rom[3962] = 12'd3962;
        rom[3963] = 12'd3963;
        rom[3964] = 12'd3964;
        rom[3965] = 12'd3965;
        rom[3966] = 12'd3966;
        rom[3967] = 12'd3967;
        rom[3968] = 12'd3968;
        rom[3969] = 12'd3969;
        rom[3970] = 12'd3970;
        rom[3971] = 12'd3971;
        rom[3972] = 12'd3972;
        rom[3973] = 12'd3973;
        rom[3974] = 12'd3974;
        rom[3975] = 12'd3975;
        rom[3976] = 12'd3976;
        rom[3977] = 12'd3977;
        rom[3978] = 12'd3978;
        rom[3979] = 12'd3979;
        rom[3980] = 12'd3980;
        rom[3981] = 12'd3981;
        rom[3982] = 12'd3982;
        rom[3983] = 12'd3983;
        rom[3984] = 12'd3984;
        rom[3985] = 12'd3985;
        rom[3986] = 12'd3986;
        rom[3987] = 12'd3987;
        rom[3988] = 12'd3988;
        rom[3989] = 12'd3989;
        rom[3990] = 12'd3990;
        rom[3991] = 12'd3991;
        rom[3992] = 12'd3992;
        rom[3993] = 12'd3993;
        rom[3994] = 12'd3994;
        rom[3995] = 12'd3995;
        rom[3996] = 12'd3996;
        rom[3997] = 12'd3997;
        rom[3998] = 12'd3998;
        rom[3999] = 12'd3999;
        rom[4000] = 12'd4000;
        rom[4001] = 12'd4001;
        rom[4002] = 12'd4002;
        rom[4003] = 12'd4003;
        rom[4004] = 12'd4004;
        rom[4005] = 12'd4005;
        rom[4006] = 12'd4006;
        rom[4007] = 12'd4007;
        rom[4008] = 12'd4008;
        rom[4009] = 12'd4009;
        rom[4010] = 12'd4010;
        rom[4011] = 12'd4011;
        rom[4012] = 12'd4012;
        rom[4013] = 12'd4013;
        rom[4014] = 12'd4014;
        rom[4015] = 12'd4015;
        rom[4016] = 12'd4016;
        rom[4017] = 12'd4017;
        rom[4018] = 12'd4018;
        rom[4019] = 12'd4019;
        rom[4020] = 12'd4020;
        rom[4021] = 12'd4021;
        rom[4022] = 12'd4022;
        rom[4023] = 12'd4023;
        rom[4024] = 12'd4024;
        rom[4025] = 12'd4025;
        rom[4026] = 12'd4026;
        rom[4027] = 12'd4027;
        rom[4028] = 12'd4028;
        rom[4029] = 12'd4029;
        rom[4030] = 12'd4030;
        rom[4031] = 12'd4031;
        rom[4032] = 12'd4032;
        rom[4033] = 12'd4033;
        rom[4034] = 12'd4034;
        rom[4035] = 12'd4035;
        rom[4036] = 12'd4036;
        rom[4037] = 12'd4037;
        rom[4038] = 12'd4038;
        rom[4039] = 12'd4039;
        rom[4040] = 12'd4040;
        rom[4041] = 12'd4041;
        rom[4042] = 12'd4042;
        rom[4043] = 12'd4043;
        rom[4044] = 12'd4044;
        rom[4045] = 12'd4045;
        rom[4046] = 12'd4046;
        rom[4047] = 12'd4047;
        rom[4048] = 12'd4048;
        rom[4049] = 12'd4049;
        rom[4050] = 12'd4050;
        rom[4051] = 12'd4051;
        rom[4052] = 12'd4052;
        rom[4053] = 12'd4053;
        rom[4054] = 12'd4054;
        rom[4055] = 12'd4055;
        rom[4056] = 12'd4056;
        rom[4057] = 12'd4057;
        rom[4058] = 12'd4058;
        rom[4059] = 12'd4059;
        rom[4060] = 12'd4060;
        rom[4061] = 12'd4061;
        rom[4062] = 12'd4062;
        rom[4063] = 12'd4063;
        rom[4064] = 12'd4064;
        rom[4065] = 12'd4065;
        rom[4066] = 12'd4066;
        rom[4067] = 12'd4067;
        rom[4068] = 12'd4068;
        rom[4069] = 12'd4069;
        rom[4070] = 12'd4070;
        rom[4071] = 12'd4071;
        rom[4072] = 12'd4072;
        rom[4073] = 12'd4073;
        rom[4074] = 12'd4074;
        rom[4075] = 12'd4075;
        rom[4076] = 12'd4076;
        rom[4077] = 12'd4077;
        rom[4078] = 12'd4078;
        rom[4079] = 12'd4079;
        rom[4080] = 12'd4080;
        rom[4081] = 12'd4081;
        rom[4082] = 12'd4082;
        rom[4083] = 12'd4083;
        rom[4084] = 12'd4084;
        rom[4085] = 12'd4085;
        rom[4086] = 12'd4086;
        rom[4087] = 12'd4087;
        rom[4088] = 12'd4088;
        rom[4089] = 12'd4089;
        rom[4090] = 12'd4090;
        rom[4091] = 12'd4091;
        rom[4092] = 12'd4092;
        rom[4093] = 12'd4093;
        rom[4094] = 12'd4094;
        rom[4095] = 12'd4095;
    end

    always @(posedge clk) begin
        if (we) rom[addr] <= di;
        dout <= rom[addr];
    end

endmodule